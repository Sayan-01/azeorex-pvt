<svg width="645" height="481" viewBox="0 0 645 481" fill="none" xmlns="http://www.w3.org/2000/svg" xmlns:xlink="http://www.w3.org/1999/xlink">
<rect width="640" height="477" transform="translate(3 4)" fill="#1E1E20"/>
<rect x="3" y="4" width="640" height="477" fill="url(#pattern0_349_17)"/>
<path d="M37.4038 447.289C35.9846 447.289 34.717 447.045 33.6009 446.556C32.4918 446.067 31.6134 445.388 30.9658 444.52C30.3251 443.645 29.9806 442.632 29.9324 441.482H33.1772C33.2186 442.109 33.4287 442.653 33.8076 443.114C34.1934 443.569 34.6963 443.921 35.3163 444.169C35.9364 444.417 36.6253 444.541 37.3831 444.541C38.2167 444.541 38.9538 444.396 39.5945 444.107C40.2421 443.817 40.7485 443.414 41.1136 442.897C41.4787 442.374 41.6613 441.771 41.6613 441.089C41.6613 440.379 41.4787 439.756 41.1136 439.219C40.7554 438.674 40.2283 438.247 39.5325 437.937C38.8436 437.627 38.01 437.472 37.0317 437.472H35.244V434.868H37.0317C37.8171 434.868 38.506 434.727 39.0985 434.444C39.6979 434.162 40.1663 433.769 40.5039 433.266C40.8415 432.757 41.0103 432.161 41.0103 431.479C41.0103 430.824 40.8621 430.256 40.5659 429.774C40.2766 429.284 39.8632 428.902 39.3259 428.626C38.7954 428.351 38.1685 428.213 37.4451 428.213C36.7562 428.213 36.112 428.341 35.5127 428.595C34.9202 428.844 34.438 429.202 34.0659 429.67C33.6939 430.132 33.4941 430.686 33.4666 431.334H30.3768C30.4112 430.19 30.7488 429.185 31.3895 428.316C32.0371 427.448 32.8913 426.77 33.9523 426.281C35.0132 425.792 36.1913 425.547 37.4864 425.547C38.8436 425.547 40.0148 425.812 40.9999 426.343C41.992 426.866 42.7567 427.566 43.294 428.44C43.8383 429.315 44.107 430.273 44.1001 431.313C44.107 432.498 43.7763 433.504 43.108 434.331C42.4467 435.157 41.5648 435.712 40.4626 435.994V436.16C41.868 436.373 42.9565 436.931 43.7281 437.834C44.5065 438.736 44.8923 439.856 44.8854 441.192C44.8923 442.357 44.5685 443.4 43.9141 444.324C43.2665 445.247 42.3812 445.974 41.2583 446.504C40.1353 447.028 38.8505 447.289 37.4038 447.289ZM49.5047 447L58.7431 428.73V428.575H48.0579V425.836H62.0499V428.668L52.8425 447H49.5047ZM73.7452 424.844L66.9249 450.183H64.1657L70.9861 424.844H73.7452ZM83.3143 447.289C82.0191 447.289 80.8548 447.041 79.8215 446.545C78.795 446.042 77.9752 445.353 77.362 444.479C76.7489 443.604 76.4216 442.605 76.3803 441.482H79.4804C79.5562 442.391 79.9592 443.139 80.6895 443.724C81.4198 444.31 82.2947 444.603 83.3143 444.603C84.1272 444.603 84.8471 444.417 85.4741 444.045C86.1079 443.666 86.6039 443.145 86.9621 442.484C87.3272 441.823 87.5098 441.068 87.5098 440.221C87.5098 439.36 87.3238 438.592 86.9518 437.917C86.5798 437.241 86.0665 436.711 85.412 436.325C84.7645 435.939 84.0204 435.743 83.1799 435.736C82.5393 435.736 81.8951 435.846 81.2475 436.067C80.5999 436.287 80.0764 436.577 79.6768 436.935L76.7523 436.501L77.9407 425.836H89.5766V428.575H80.5965L79.9248 434.496H80.0488C80.4622 434.097 81.0098 433.762 81.6919 433.494C82.3808 433.225 83.1179 433.091 83.9033 433.091C85.1916 433.091 86.3386 433.397 87.3445 434.01C88.3572 434.624 89.1529 435.461 89.7316 436.522C90.3172 437.576 90.6065 438.788 90.5996 440.159C90.6065 441.53 90.2965 442.753 89.6696 443.828C89.0496 444.902 88.1884 445.75 87.0861 446.37C85.9907 446.983 84.7335 447.289 83.3143 447.289ZM93.9297 442.866V440.283L103.075 425.836H105.111V429.639H103.819L97.2778 439.994V440.159H109.813V442.866H93.9297ZM103.964 447V442.081L103.984 440.903V425.836H107.012V447H103.964ZM121.157 447V431.127H124.143V433.649H124.308C124.598 432.794 125.108 432.123 125.838 431.634C126.575 431.138 127.409 430.89 128.339 430.89C128.532 430.89 128.759 430.896 129.021 430.91C129.289 430.924 129.5 430.941 129.651 430.962V433.917C129.527 433.883 129.307 433.845 128.99 433.804C128.673 433.756 128.356 433.731 128.039 433.731C127.309 433.731 126.658 433.886 126.086 434.196C125.521 434.5 125.073 434.923 124.743 435.467C124.412 436.005 124.246 436.618 124.246 437.307V447H121.157ZM138.598 447.32C137.034 447.32 135.687 446.986 134.557 446.318C133.434 445.643 132.566 444.696 131.953 443.476C131.347 442.25 131.044 440.813 131.044 439.167C131.044 437.541 131.347 436.108 131.953 434.868C132.566 433.628 133.42 432.66 134.516 431.964C135.618 431.269 136.906 430.921 138.381 430.921C139.276 430.921 140.144 431.069 140.985 431.365C141.825 431.661 142.58 432.126 143.248 432.76C143.916 433.394 144.443 434.217 144.829 435.23C145.215 436.236 145.408 437.458 145.408 438.898V439.994H132.79V437.679H142.38C142.38 436.866 142.214 436.146 141.884 435.519C141.553 434.885 141.088 434.386 140.489 434.021C139.896 433.656 139.2 433.473 138.401 433.473C137.533 433.473 136.775 433.687 136.128 434.114C135.487 434.534 134.991 435.085 134.64 435.767C134.295 436.442 134.123 437.176 134.123 437.968V439.777C134.123 440.838 134.309 441.74 134.681 442.484C135.06 443.228 135.587 443.797 136.262 444.189C136.937 444.575 137.726 444.768 138.629 444.768C139.214 444.768 139.748 444.685 140.23 444.52C140.713 444.348 141.129 444.093 141.481 443.755C141.832 443.418 142.101 443.001 142.287 442.505L145.211 443.032C144.977 443.893 144.557 444.647 143.95 445.295C143.351 445.936 142.597 446.435 141.687 446.793C140.785 447.145 139.755 447.32 138.598 447.32ZM160.73 435.002L157.93 435.498C157.812 435.14 157.626 434.799 157.372 434.475C157.123 434.152 156.786 433.886 156.359 433.68C155.932 433.473 155.398 433.37 154.757 433.37C153.882 433.37 153.152 433.566 152.566 433.959C151.981 434.345 151.688 434.844 151.688 435.457C151.688 435.988 151.884 436.415 152.277 436.739C152.67 437.062 153.303 437.328 154.178 437.534L156.7 438.113C158.16 438.45 159.249 438.971 159.965 439.673C160.682 440.376 161.04 441.289 161.04 442.412C161.04 443.362 160.764 444.21 160.213 444.954C159.669 445.691 158.908 446.27 157.93 446.69C156.958 447.11 155.832 447.32 154.55 447.32C152.773 447.32 151.323 446.941 150.2 446.184C149.077 445.419 148.388 444.334 148.133 442.928L151.12 442.474C151.306 443.252 151.688 443.841 152.267 444.241C152.845 444.634 153.6 444.83 154.53 444.83C155.542 444.83 156.352 444.62 156.958 444.2C157.564 443.772 157.868 443.252 157.868 442.639C157.868 442.143 157.682 441.726 157.31 441.389C156.944 441.051 156.383 440.796 155.625 440.624L152.938 440.035C151.457 439.697 150.362 439.16 149.652 438.423C148.949 437.686 148.598 436.752 148.598 435.622C148.598 434.686 148.86 433.866 149.383 433.163C149.907 432.46 150.63 431.913 151.554 431.52C152.477 431.12 153.534 430.921 154.726 430.921C156.441 430.921 157.792 431.293 158.777 432.037C159.762 432.774 160.413 433.762 160.73 435.002ZM171.123 447.32C169.635 447.32 168.337 446.979 167.227 446.297C166.118 445.615 165.257 444.661 164.644 443.435C164.031 442.209 163.724 440.776 163.724 439.136C163.724 437.489 164.031 436.05 164.644 434.816C165.257 433.583 166.118 432.626 167.227 431.944C168.337 431.262 169.635 430.921 171.123 430.921C172.611 430.921 173.91 431.262 175.019 431.944C176.128 432.626 176.989 433.583 177.603 434.816C178.216 436.05 178.522 437.489 178.522 439.136C178.522 440.776 178.216 442.209 177.603 443.435C176.989 444.661 176.128 445.615 175.019 446.297C173.91 446.979 172.611 447.32 171.123 447.32ZM171.134 444.727C172.098 444.727 172.897 444.472 173.531 443.962C174.165 443.452 174.633 442.773 174.936 441.926C175.246 441.079 175.401 440.145 175.401 439.126C175.401 438.113 175.246 437.183 174.936 436.336C174.633 435.481 174.165 434.796 173.531 434.279C172.897 433.762 172.098 433.504 171.134 433.504C170.162 433.504 169.356 433.762 168.715 434.279C168.082 434.796 167.61 435.481 167.3 436.336C166.997 437.183 166.845 438.113 166.845 439.126C166.845 440.145 166.997 441.079 167.3 441.926C167.61 442.773 168.082 443.452 168.715 443.962C169.356 444.472 170.162 444.727 171.134 444.727ZM185.061 425.836V447H181.971V425.836H185.061ZM202.796 431.127L197.04 447H193.734L187.967 431.127H191.284L195.304 443.342H195.47L199.479 431.127H202.796ZM212.001 447.32C210.437 447.32 209.091 446.986 207.961 446.318C206.838 445.643 205.97 444.696 205.357 443.476C204.75 442.25 204.447 440.813 204.447 439.167C204.447 437.541 204.75 436.108 205.357 434.868C205.97 433.628 206.824 432.66 207.919 431.964C209.022 431.269 210.31 430.921 211.784 430.921C212.68 430.921 213.548 431.069 214.388 431.365C215.229 431.661 215.983 432.126 216.651 432.76C217.32 433.394 217.847 434.217 218.232 435.23C218.618 436.236 218.811 437.458 218.811 438.898V439.994H206.194V437.679H215.783C215.783 436.866 215.618 436.146 215.287 435.519C214.957 434.885 214.492 434.386 213.892 434.021C213.3 433.656 212.604 433.473 211.805 433.473C210.937 433.473 210.179 433.687 209.531 434.114C208.891 434.534 208.395 435.085 208.043 435.767C207.699 436.442 207.527 437.176 207.527 437.968V439.777C207.527 440.838 207.713 441.74 208.085 442.484C208.464 443.228 208.991 443.797 209.666 444.189C210.341 444.575 211.13 444.768 212.032 444.768C212.618 444.768 213.152 444.685 213.634 444.52C214.116 444.348 214.533 444.093 214.884 443.755C215.236 443.418 215.504 443.001 215.69 442.505L218.615 443.032C218.381 443.893 217.96 444.647 217.354 445.295C216.755 445.936 216 446.435 215.091 446.793C214.189 447.145 213.159 447.32 212.001 447.32ZM228.181 447.31C226.9 447.31 225.756 446.983 224.751 446.328C223.752 445.667 222.966 444.727 222.394 443.507C221.829 442.281 221.547 440.81 221.547 439.095C221.547 437.379 221.833 435.912 222.405 434.692C222.983 433.473 223.776 432.54 224.782 431.892C225.787 431.244 226.928 430.921 228.202 430.921C229.187 430.921 229.979 431.086 230.579 431.417C231.185 431.74 231.654 432.119 231.984 432.553C232.322 432.987 232.584 433.37 232.77 433.7H232.956V425.836H236.045V447H233.028V444.53H232.77C232.584 444.868 232.315 445.254 231.964 445.688C231.619 446.122 231.144 446.501 230.537 446.824C229.931 447.148 229.146 447.31 228.181 447.31ZM228.863 444.675C229.752 444.675 230.503 444.441 231.116 443.972C231.736 443.497 232.205 442.839 232.522 441.998C232.845 441.158 233.007 440.18 233.007 439.064C233.007 437.961 232.849 436.997 232.532 436.17C232.215 435.343 231.75 434.699 231.137 434.238C230.524 433.776 229.766 433.545 228.863 433.545C227.933 433.545 227.158 433.787 226.538 434.269C225.918 434.751 225.45 435.409 225.133 436.243C224.823 437.076 224.668 438.016 224.668 439.064C224.668 440.125 224.826 441.079 225.143 441.926C225.46 442.773 225.929 443.445 226.549 443.941C227.176 444.43 227.947 444.675 228.863 444.675Z" fill="#6D6D6F"/>
<path d="M48.0012 367.764H51.8212V384.362C51.8212 386.128 51.4063 387.693 50.5766 389.057C49.7469 390.412 48.5804 391.48 47.077 392.261C45.5737 393.033 43.8116 393.419 41.7907 393.419C39.778 393.419 38.02 393.033 36.5167 392.261C35.0134 391.48 33.8468 390.412 33.0171 389.057C32.1874 387.693 31.7725 386.128 31.7725 384.362V367.764H35.5802V384.054C35.5802 385.196 35.8307 386.21 36.3319 387.098C36.8412 387.985 37.56 388.683 38.4883 389.192C39.4166 389.693 40.5174 389.944 41.7907 389.944C43.0722 389.944 44.1771 389.693 45.1054 389.192C46.0419 388.683 46.7566 387.985 47.2495 387.098C47.7507 386.21 48.0012 385.196 48.0012 384.054V367.764ZM60.7457 381.762V393H57.0613V374.073H60.5978V377.153H60.832C61.2673 376.151 61.9492 375.346 62.8775 374.738C63.814 374.13 64.9928 373.826 66.414 373.826C67.7038 373.826 68.8333 374.097 69.8027 374.64C70.7721 375.174 71.5237 375.97 72.0577 377.03C72.5917 378.09 72.8587 379.4 72.8587 380.961V393H69.1742V381.405C69.1742 380.033 68.8169 378.961 68.1022 378.188C67.3875 377.408 66.4058 377.018 65.1571 377.018C64.3028 377.018 63.5429 377.203 62.8775 377.572C62.2203 377.942 61.6986 378.484 61.3125 379.199C60.9346 379.905 60.7457 380.76 60.7457 381.762ZM86.6351 374.073V377.03H76.2966V374.073H86.6351ZM79.0692 369.538H82.7536V387.443C82.7536 388.157 82.8604 388.695 83.074 389.057C83.2875 389.41 83.5628 389.652 83.8996 389.784C84.2446 389.907 84.6184 389.969 85.0209 389.969C85.3166 389.969 85.5754 389.948 85.7972 389.907C86.019 389.866 86.1915 389.833 86.3148 389.808L86.9802 392.852C86.7666 392.934 86.4626 393.016 86.0683 393.099C85.674 393.189 85.1811 393.238 84.5896 393.246C83.6203 393.263 82.7166 393.09 81.8787 392.729C81.0408 392.367 80.363 391.809 79.8455 391.053C79.3279 390.297 79.0692 389.348 79.0692 388.207V369.538ZM90.7108 393V374.073H94.3952V393H90.7108ZM92.5715 371.152C91.9307 371.152 91.3803 370.939 90.9203 370.512C90.4685 370.076 90.2425 369.559 90.2425 368.959C90.2425 368.351 90.4685 367.833 90.9203 367.406C91.3803 366.971 91.9307 366.753 92.5715 366.753C93.2123 366.753 93.7585 366.971 94.2104 367.406C94.6704 367.833 94.9004 368.351 94.9004 368.959C94.9004 369.559 94.6704 370.076 94.2104 370.512C93.7585 370.939 93.2123 371.152 92.5715 371.152ZM108.187 374.073V377.03H97.8486V374.073H108.187ZM100.621 369.538H104.306V387.443C104.306 388.157 104.412 388.695 104.626 389.057C104.84 389.41 105.115 389.652 105.452 389.784C105.797 389.907 106.17 389.969 106.573 389.969C106.869 389.969 107.127 389.948 107.349 389.907C107.571 389.866 107.743 389.833 107.867 389.808L108.532 392.852C108.319 392.934 108.015 393.016 107.62 393.099C107.226 393.189 106.733 393.238 106.142 393.246C105.172 393.263 104.269 393.09 103.431 392.729C102.593 392.367 101.915 391.809 101.397 391.053C100.88 390.297 100.621 389.348 100.621 388.207V369.538ZM116.354 367.764V393H112.669V367.764H116.354ZM129.468 393.382C127.603 393.382 125.997 392.984 124.65 392.187C123.311 391.382 122.276 390.252 121.545 388.798C120.822 387.336 120.46 385.623 120.46 383.66C120.46 381.721 120.822 380.012 121.545 378.533C122.276 377.055 123.294 375.901 124.601 375.071C125.915 374.241 127.451 373.826 129.209 373.826C130.277 373.826 131.312 374.003 132.314 374.356C133.317 374.709 134.216 375.264 135.013 376.02C135.81 376.775 136.438 377.757 136.898 378.965C137.358 380.164 137.588 381.622 137.588 383.339V384.645H122.543V381.885H133.978C133.978 380.916 133.781 380.057 133.387 379.31C132.992 378.554 132.438 377.958 131.723 377.523C131.016 377.088 130.187 376.87 129.234 376.87C128.199 376.87 127.295 377.125 126.523 377.634C125.759 378.135 125.167 378.792 124.748 379.606C124.338 380.411 124.132 381.285 124.132 382.23V384.387C124.132 385.652 124.354 386.728 124.798 387.615C125.25 388.502 125.878 389.18 126.683 389.648C127.488 390.108 128.429 390.338 129.505 390.338C130.203 390.338 130.84 390.24 131.415 390.043C131.99 389.837 132.487 389.533 132.906 389.131C133.325 388.728 133.645 388.231 133.867 387.64L137.354 388.268C137.075 389.295 136.574 390.195 135.851 390.967C135.136 391.731 134.237 392.326 133.152 392.754C132.076 393.173 130.848 393.382 129.468 393.382ZM148.762 393.37C147.234 393.37 145.87 392.979 144.671 392.199C143.48 391.41 142.543 390.289 141.861 388.835C141.188 387.373 140.851 385.619 140.851 383.573C140.851 381.528 141.192 379.778 141.874 378.324C142.564 376.87 143.508 375.757 144.708 374.985C145.907 374.212 147.267 373.826 148.786 373.826C149.961 373.826 150.906 374.023 151.621 374.418C152.344 374.804 152.902 375.256 153.296 375.773C153.699 376.291 154.011 376.747 154.233 377.141H154.455V367.764H158.139V393H154.541V390.055H154.233C154.011 390.457 153.691 390.918 153.272 391.435C152.861 391.953 152.294 392.404 151.571 392.791C150.848 393.177 149.912 393.37 148.762 393.37ZM149.575 390.227C150.635 390.227 151.53 389.948 152.261 389.39C153.001 388.823 153.559 388.038 153.937 387.036C154.323 386.034 154.516 384.867 154.516 383.536C154.516 382.222 154.327 381.072 153.95 380.086C153.572 379.1 153.017 378.332 152.286 377.782C151.555 377.231 150.651 376.956 149.575 376.956C148.466 376.956 147.542 377.244 146.803 377.819C146.063 378.394 145.505 379.178 145.127 380.172C144.757 381.166 144.572 382.288 144.572 383.536C144.572 384.801 144.761 385.939 145.139 386.95C145.517 387.96 146.076 388.761 146.815 389.353C147.562 389.936 148.483 390.227 149.575 390.227ZM172.877 393V367.764H181.872C183.836 367.764 185.462 368.121 186.752 368.836C188.042 369.55 189.007 370.528 189.648 371.768C190.288 373.001 190.609 374.389 190.609 375.933C190.609 377.486 190.284 378.883 189.635 380.123C188.995 381.355 188.025 382.333 186.727 383.056C185.438 383.77 183.815 384.128 181.86 384.128H175.674V380.899H181.515C182.755 380.899 183.762 380.686 184.534 380.259C185.306 379.823 185.873 379.232 186.234 378.484C186.596 377.737 186.777 376.886 186.777 375.933C186.777 374.98 186.596 374.134 186.234 373.395C185.873 372.656 185.302 372.076 184.522 371.658C183.749 371.239 182.731 371.029 181.466 371.029H176.684V393H172.877ZM194.777 393V374.073H198.338V377.079H198.535C198.88 376.061 199.488 375.26 200.359 374.677C201.238 374.085 202.232 373.789 203.341 373.789C203.571 373.789 203.842 373.798 204.154 373.814C204.475 373.83 204.725 373.851 204.906 373.876V377.4C204.758 377.359 204.495 377.314 204.117 377.264C203.739 377.207 203.362 377.178 202.984 377.178C202.113 377.178 201.337 377.363 200.655 377.732C199.981 378.094 199.447 378.599 199.053 379.248C198.658 379.889 198.461 380.62 198.461 381.442V393H194.777ZM215.389 393.382C213.615 393.382 212.066 392.975 210.744 392.162C209.421 391.349 208.394 390.211 207.663 388.749C206.932 387.286 206.566 385.578 206.566 383.623C206.566 381.659 206.932 379.942 207.663 378.472C208.394 377.001 209.421 375.859 210.744 375.046C212.066 374.233 213.615 373.826 215.389 373.826C217.164 373.826 218.712 374.233 220.035 375.046C221.357 375.859 222.384 377.001 223.115 378.472C223.847 379.942 224.212 381.659 224.212 383.623C224.212 385.578 223.847 387.286 223.115 388.749C222.384 390.211 221.357 391.349 220.035 392.162C218.712 392.975 217.164 393.382 215.389 393.382ZM215.402 390.289C216.552 390.289 217.505 389.985 218.26 389.377C219.016 388.769 219.575 387.96 219.936 386.95C220.306 385.939 220.491 384.826 220.491 383.61C220.491 382.403 220.306 381.294 219.936 380.283C219.575 379.265 219.016 378.447 218.26 377.831C217.505 377.215 216.552 376.907 215.402 376.907C214.243 376.907 213.282 377.215 212.518 377.831C211.762 378.447 211.2 379.265 210.83 380.283C210.469 381.294 210.288 382.403 210.288 383.61C210.288 384.826 210.469 385.939 210.83 386.95C211.2 387.96 211.762 388.769 212.518 389.377C213.282 389.985 214.243 390.289 215.402 390.289ZM228.325 374.073H232.009V394.232C232.009 395.497 231.779 396.565 231.319 397.436C230.867 398.307 230.194 398.968 229.298 399.42C228.411 399.872 227.314 400.098 226.008 400.098C225.877 400.098 225.753 400.098 225.638 400.098C225.515 400.098 225.388 400.094 225.256 400.085V396.919C225.371 396.919 225.474 396.919 225.565 396.919C225.647 396.919 225.741 396.919 225.848 396.919C226.719 396.919 227.347 396.684 227.733 396.216C228.128 395.756 228.325 395.087 228.325 394.208V374.073ZM230.148 371.152C229.508 371.152 228.957 370.939 228.497 370.512C228.045 370.076 227.82 369.559 227.82 368.959C227.82 368.351 228.045 367.833 228.497 367.406C228.957 366.971 229.508 366.753 230.148 366.753C230.789 366.753 231.336 366.971 231.787 367.406C232.247 367.833 232.477 368.351 232.477 368.959C232.477 369.559 232.247 370.076 231.787 370.512C231.336 370.939 230.789 371.152 230.148 371.152ZM245.123 393.382C243.259 393.382 241.653 392.984 240.305 392.187C238.966 391.382 237.931 390.252 237.2 388.798C236.477 387.336 236.116 385.623 236.116 383.66C236.116 381.721 236.477 380.012 237.2 378.533C237.931 377.055 238.95 375.901 240.256 375.071C241.57 374.241 243.107 373.826 244.865 373.826C245.933 373.826 246.968 374.003 247.97 374.356C248.972 374.709 249.872 375.264 250.668 376.02C251.465 376.775 252.094 377.757 252.554 378.965C253.014 380.164 253.244 381.622 253.244 383.339V384.645H238.198V381.885H249.633C249.633 380.916 249.436 380.057 249.042 379.31C248.648 378.554 248.093 377.958 247.378 377.523C246.672 377.088 245.842 376.87 244.889 376.87C243.854 376.87 242.95 377.125 242.178 377.634C241.414 378.135 240.823 378.792 240.404 379.606C239.993 380.411 239.788 381.285 239.788 382.23V384.387C239.788 385.652 240.01 386.728 240.453 387.615C240.905 388.502 241.533 389.18 242.338 389.648C243.144 390.108 244.084 390.338 245.16 390.338C245.859 390.338 246.495 390.24 247.07 390.043C247.645 389.837 248.142 389.533 248.561 389.131C248.98 388.728 249.301 388.231 249.522 387.64L253.01 388.268C252.73 389.295 252.229 390.195 251.506 390.967C250.792 391.731 249.892 392.326 248.808 392.754C247.732 393.173 246.503 393.382 245.123 393.382ZM265.304 393.382C263.472 393.382 261.895 392.967 260.573 392.137C259.258 391.3 258.248 390.145 257.541 388.675C256.835 387.204 256.482 385.52 256.482 383.623C256.482 381.7 256.843 380.004 257.566 378.533C258.289 377.055 259.307 375.901 260.622 375.071C261.936 374.241 263.485 373.826 265.267 373.826C266.705 373.826 267.987 374.093 269.112 374.627C270.237 375.153 271.145 375.892 271.835 376.845C272.534 377.798 272.948 378.911 273.08 380.185H269.494C269.297 379.297 268.845 378.533 268.139 377.893C267.44 377.252 266.504 376.932 265.329 376.932C264.302 376.932 263.403 377.203 262.63 377.745C261.866 378.279 261.271 379.043 260.844 380.037C260.417 381.023 260.203 382.189 260.203 383.536C260.203 384.916 260.412 386.108 260.831 387.11C261.25 388.112 261.842 388.888 262.606 389.439C263.378 389.989 264.286 390.264 265.329 390.264C266.027 390.264 266.66 390.137 267.227 389.882C267.802 389.62 268.282 389.246 268.668 388.761C269.063 388.276 269.338 387.693 269.494 387.011H273.08C272.948 388.235 272.55 389.328 271.885 390.289C271.219 391.25 270.328 392.006 269.211 392.556C268.102 393.107 266.8 393.382 265.304 393.382ZM285.855 374.073V377.03H275.517V374.073H285.855ZM278.289 369.538H281.974V387.443C281.974 388.157 282.08 388.695 282.294 389.057C282.508 389.41 282.783 389.652 283.12 389.784C283.465 389.907 283.838 389.969 284.241 389.969C284.537 389.969 284.795 389.948 285.017 389.907C285.239 389.866 285.412 389.833 285.535 389.808L286.2 392.852C285.987 392.934 285.683 393.016 285.288 393.099C284.894 393.189 284.401 393.238 283.81 393.246C282.84 393.263 281.937 393.09 281.099 392.729C280.261 392.367 279.583 391.809 279.066 391.053C278.548 390.297 278.289 389.348 278.289 388.207V369.538Z" fill="#CDCDCF"/>
<rect width="645" height="337" fill="url(#pattern1_349_17)"/>
<path d="M295.252 186V163.164H303.816C305.57 163.164 307.042 163.491 308.232 164.145C309.429 164.799 310.332 165.699 310.941 166.843C311.558 167.981 311.867 169.274 311.867 170.724C311.867 172.188 311.558 173.489 310.941 174.626C310.324 175.764 309.414 176.66 308.209 177.314C307.005 177.96 305.522 178.284 303.76 178.284H298.085V174.883H303.203C304.229 174.883 305.069 174.704 305.723 174.348C306.377 173.991 306.86 173.5 307.172 172.876C307.492 172.251 307.652 171.534 307.652 170.724C307.652 169.913 307.492 169.2 307.172 168.583C306.86 167.966 306.373 167.486 305.712 167.144C305.057 166.795 304.214 166.62 303.18 166.62H299.389V186H295.252ZM315.46 186V163.164H324.024C325.778 163.164 327.25 163.468 328.439 164.078C329.636 164.688 330.539 165.542 331.149 166.643C331.766 167.735 332.074 169.01 332.074 170.467C332.074 171.932 331.762 173.203 331.138 174.281C330.521 175.351 329.61 176.18 328.406 176.767C327.202 177.347 325.722 177.637 323.968 177.637H317.869V174.203H323.41C324.436 174.203 325.276 174.061 325.93 173.779C326.585 173.489 327.068 173.069 327.38 172.519C327.7 171.961 327.859 171.278 327.859 170.467C327.859 169.657 327.7 168.966 327.38 168.393C327.06 167.813 326.573 167.375 325.919 167.077C325.265 166.773 324.421 166.62 323.388 166.62H319.597V186H315.46ZM327.257 175.652L332.911 186H328.294L322.741 175.652H327.257ZM344.892 163.164H348.995V179.22C348.988 180.692 348.676 181.96 348.059 183.023C347.442 184.078 346.579 184.892 345.472 185.465C344.372 186.03 343.089 186.312 341.625 186.312C340.287 186.312 339.083 186.074 338.012 185.599C336.949 185.115 336.105 184.402 335.481 183.458C334.856 182.514 334.544 181.339 334.544 179.934H338.659C338.666 180.551 338.8 181.083 339.06 181.529C339.328 181.975 339.696 182.317 340.164 182.554C340.632 182.792 341.171 182.911 341.781 182.911C342.443 182.911 343.004 182.774 343.465 182.499C343.926 182.216 344.275 181.8 344.513 181.25C344.758 180.7 344.885 180.023 344.892 179.22V163.164Z" fill="#B2B5B4"/>
<defs>
<pattern id="pattern0_349_17" patternContentUnits="objectBoundingBox" width="1" height="1">
<use xlink:href="#image0_349_17" transform="matrix(0.0015625 0 0 0.00209644 -0.0125 -0.00838575)"/>
</pattern>
<pattern id="pattern1_349_17" patternContentUnits="objectBoundingBox" width="1" height="1">
<use xlink:href="#image1_349_17" transform="scale(0.00155039 0.00296736)"/>
</pattern>
<image id="image0_349_17" width="655" height="490" preserveAspectRatio="none" xlink:href="data:image/png;base64,iVBORw0KGgoAAAANSUhEUgAAAo8AAAHqCAYAAABlQaQPAAAWy0lEQVR4nO3dW1Mi2baA0bkSvJRdt+69++XsiI7z/39bxz5d5RWEXOcBoRARJoiaiWN0VFS1CiSZKJ9r5aX89df/1lhR65MPAQDwwZRSnnyseYflAACgp8QjAABp4hEAgDTxCABAmngEACBNPAIAkCYeAQBIE48AAKSJRwAA0sQjAABp4hEAgDTxCABAmngEACBNPAIAkCYeAQBIE48AAKSJRwAA0sQjAABp4hEAgDTxCABAmngEAGCtUsqTjw3fYTkAAOiJ1YA08ggAQJp4BAAgzbQ1AABr1VoX/55PXxt5BAAgTTwCAJAmHgEASLPPIwAAay3v8zhn5BEAgDTxCABAmngEACBNPAIAkCYeAQBIE48AAKSJRwAA0sQjAABp4hEAgDTxCABAmngEACBNPAIAkCYeAQBIE48AAKSJRwAA0sQjAABp4hEAgDTxCABAmngEACBt+N4LAABAN5VSnnzMyCMAAGniEQCANPEIAECaeAQAIE08AgCQJh4BAEgTjwAApIlHAADSxCMAAGniEQCANPEIAECaeAQAIE08AgCQJh4BAEgTjwAApIlHAADSxCMAAGniEQCANPEIAECaeAQAIE08AgCQJh4BAEgTjwAApIlHAADSxCMAAGniEQCANPEIAECaeAQAIE08AgCQJh4BAEgTjwAApIlHAADSxCMAAGniEQCANPEIAECaeAQAIE08AgCQJh4BAEgTjwAApIlHAADSxCMAAGniEQCANPEIAECaeAQAIE08AgCQJh4BAEgTjwAApIlHAADSxCMAAGniEQCANPEIAECaeAQAIE08AgCQJh4BAEgTjwAApIlHAADSxCMAAGniEQCANPEIAECaeAQAIE08AgCQJh4BAEgTjwAApIlHAADSxCMAAGniEQCANPEIAECaeAQAIE08AgCQJh4BAEgTjwAApIlHAADSxCMAAGniEQCANPEIAECaeAQAIE08AgCQJh4BAEgTjwAApIlHAADSxCMAAGniEQCANPEIAECaeAQAIE08AgCQJh4BAEgTjwAApIlHAADSxCMAAGniEQCANPEIAECaeAQAIE08AgCQJh4BAEgTjwAApIlHAADSxCMAAGniEQCANPEIAECaeAQAIE08AgCQJh4BAEgTjwAApIlHAADSxCMAAGniEQCANPEIAECaeAQAIE08AgCQJh4BAEgTjwAApIlHAADSxCMAAGniEQCANPEIAECaeAQAIE08AgCQJh4BAEgTjwAApIlHAADSxCMAAGniEQCANPEIAECaeAQAIE08AgCQJh4BAEgTjwAApIlHAADSxCMAAGniEQCANPEIAECaeAQAIE08AgCQJh4BAEgTjwAApIlHAADSxCMAAGniEQCANPEIAECaeAQAIE08AgCQJh4BAEgTjwAApIlHAADSxCMAAGniEQCANPEIAECaeAQAIE08AgCQJh4BAEgTjwAApIlHAADSxCMAAGniEQCANPEIAECaeAQAIE08AgCQJh4BAEgTjwAApIlHAADSxCMAAGniEQCANPEIAECaeAQAIE08AgCQJh4BAEgTjwAApIlHAADSxCMAAGniEQCANPEIAECaeAQAIE08AgCQJh4BAEgTjwAApIlHAADSxCMAAGniEQCANPEIAECaeAQAIE08AgCQJh4BAEgTjwAApIlHAADSxCMAAGniEQCANPEIAECaeAQAIE08AgCQJh4BAEgTjwAApIlHAADSxCMAAGniEQCANPEIAECaeAQAIE08AgCQJh4BAEgTjwAApIlHAADSxCMAAGniEQCANPEIAECaeAQAIE08AgCQJh4BAEgTjwAApIlHAADSxCMAAGniEQCANPEIAECaeAQAIE08AgCQJh4BAEgTjwAApIlHAADSxCMAAGniEQCANPEIAECaeAQAIE08AgCQJh4BAEgTjwAApIlHAADSxCMAAGniEQCANPEIAECaeAQAIE08AgCQJh4BAEgTjwAApIlHAADSxCMAAGniEQCANPEIAECaeAQAIE08AgCQJh4BAEgTjwAApIlHAADSxCMAAGniEQCANPEIAECaeAQAIE08AgCQJh4BAEgTjwAApIlHAADSxCMAAGniEQCANPEIAECaeAQAIE08AgCQJh4BAEgTjwAApIlHAADSxCMAAGniEQCANPEIAECaeAQAIE08AgCQJh4BAEgTjwAApIlHAADSxCMAAGniEQCANPEIAECaeAQAIE08AgCQJh4BAEgTjwAApIlHAADSxCMAAGniEQCANPEIAECaeAQAIE08AgCQJh4BAEgTjwAApIlHAADSxCMAAGniEQCANPEIAECaeAQAIE08AgCQJh4BAEgTjwAApA3XfbCUEqWUmE6n8Z//+U9cXl3G/f19lFKiKU97s0aNWuuzD1JKiRJl74Vsa7v3bfts0zrdppTN63vbfW+7/bFafX0vv/ZKlMV6WX7Nz/9eXWfPfbwpzeJ+l7fDsazz1ddWl5/Xpu29zku+J1e9dL0cclkOad3rfdmx/DzPrv9t6yP1WFveY7fZ5zHf87H3aYpj/pn6lpqmifOz8xiNR3F1eRWDwWDt96yRRwAA0taOPO6qRImNA4t19psEu3nN35r8Rpbz3Hqa/9Zboz7/NSsfX/4+KaVErY9v29WRpG2ePM8ev7Y2LnuNzT/ndvTS7d2X9dzX1/U2+67/fdfHS7b3e77WDjpa//AzdN1M5rqfqbyeg8RjxPqNOVcf/oO+2bi7RYnY5WW9/EOtRDma74lj+oG98edYqTttb2aO5XV+KPusjxIv3PUr9t9V4D0fe83CPLssx/QztQ9MWwMAkCYeAQBIS09bL44s3WNY2FAyfbHL/jm7vq7b2m6c/jmWqd8+ec3tvY3tTVaN99tl4j0fe9Wx7j/bRzvv8ygEOWav/fr2/dMttgd98Z6v1S59n3RpWT4y09YAAKSJRwAA0sQjAABp4hEAgDTxCABAmngEACBNPAIAkCYeAQBIE48AAKSJRwAA0sQjAABp4hEAgDTxCABAmngEACBNPAIAkCYeAQBIE48AAKQN33sBXqrW+uznSilvuCTbbVqeTc9jF9vup2vrBADol97H4zarMfUR46nWunje8/XxUdbDrlH+UdYLAOzLtPUHcaiRTQDgY+v9yGOJ9SNFNcTSnNE0AOBQOhWPz4Xglhs9UaOGdgQAOLxOxeM8BPeKyAemZ/s10pjZXi95Pk9uW41Kv6fX3t4AvL5uxeMBvSRA6acSJWrUJ9u+1rr4+OqBQwDAbo42HnmZZ0d/1ozclShrdx/Y5jUCbjUcSylrRx9ni1yire3Bl+GY7PJLmBFdgI+hk/G4bvSIbiilLAJyEX8l9t7HtJRyuIhM7vZQSpmNUhp9fFZTmt1i0KoE+DA6GY90V436KPj6vH/aR4nI7DZa3qZGEQF4jnhkvQ3t0Ebb2eDadcS6q88DALpKPPKhDZpBRMwi0v6PCYs9FX7t57rPKKXdUgD6Szzy5pYvl9glgmYHZfmfJWp5CMhkR24MzpVPdfG1AvCRiUcOrm9TwfOQsa/ffub7wM5PlbTxa5OBbjsAdJd45CjsPWq4Osq1PIqWvM2HsOU5Z9a/IAQ4DuKRg+nbiOMyp4c6jNUp5nkw1pq/ZKjIBOi2o4/H5SDo0pvScmhtu+rJ8omu+xxob2F5Gz8Xg6vrcO1Jzx9/wa9/lMePcPQO8XKr+59IHoDuOcp4XBcNmZGlJ6MmLwi1Go9HWjadDHvT4yxH4zEdOPBqz6cu/3N2BPX8iOppO3168uuHq82k77qW5f/jwA560ngAXsVRxuM660Y+1o1E7vrGte3rVx93nzfGtZG1dDWV5VCdf+1zYZY5ufcuy9j1N/qmNI9Pfv3w772nqXeIzV57jc26Zb3ZbQCgHzoVj4e4asmzU5Vr3g23vVk9ufxeWT8N/tx0+Ku/GS6fc2/N555Mxy6t163Rt+7TPXlvr7WuX9a65fNHKjOVv+pQo8KPvl+2vObacJ5NgD7oRDw+2f+vbn4j2fm6u8vnpHvJtNhzN9t0dweOlMyb+uKUMy8ZPepjXG3t4QMNpy1W7duPui7v/7pYnH1+EVh33w8b/eC/9Ow4038Ml74EOGadiMc+mE8Pd+mgm9WR0Kxn9zfcNJLZdR3aLK9l3+2y6xR95per7AFci++XXX7XE40AnXaU8bj6htXLGHoPO6ym1XXahX0ft56fsc9e8hJeOYgo+3iZ75uN+85GffS6mO8u0ESTWwYAOqlz8XjI0HPuvu5a3i6ZK5Ns85Lblyjp3RlKlDffN28xnfyCEbld1898m+w92lln4bj2NEjP3GV5+M81xgG6rXPx2NZ265tkp6aO6YRdQmf+tcuvo+zI6bsc1NGz33+Ww3F1f+Zt28n3NkD3dXL+aJerUfy6Ufy6jfefN7fuQI6takSp719GG8+zucPRwq+irPz9xurSfxlt20ats/Nrrltfta0xrdOY1umhFxWAN9K5kce5+ZvV1tPpJL+Oblidrv6odnruPVlN03aaC2xXnAHotc7GY0T8GkFMnlz4EPvO8TKpUwnNN+hH2VRHHknTdrpbDNdfB9M4shqgf7odj/H4Mn9rTw/ivadXXnO0MTutvBwsm05ZtM99r7V0VZp9Rl67+AtRW9tH62mfg1xW16mQBOiHzsfjOosRC+81vdCnEabnlvWgyz+/YlHPrDvA6KX7ga67dCQA3dareOzqm0tfwuiQurotXsPqZR2fXBFpzb836eJI4j4OFY6rPuL3E0Cf9CoeX9v8HHPH+uZVSonpdHrQ53es6ypjeZRyfo7CYwlDAHhOJ+Lx4AGydHWMUkpq37LFUdv7jCQdeFr2tYLsJeH4Ksu0fM3xF+6D8NYR++T60i+9lvgr2mfd7HKJwkPdHwD90Il4XLX3G9f8QzU/NZg+UfSGy7W9drgc4iATb96HsxhtXBeQrPWRR6gBjk0n4zGtZ+/VfQm4dRH0kS4b+ZYH+HR9XRyaiATov37H47IdpkCfvIG9VdOV3QLyxVO5j1fKweL1oMt1gPs7pOdGD19rGQ95v4cOfABYp5PxuMvoRInHl8Xb9coVb3qli6Xz/WW8ZJTmyfPa8bG33v+RjiA9Cduy+f9fWzbisvv2ZnUp6AHolk7GI/Ag0Y5CD4C3JB7hHS2O0t61/zYcwAUAr0k8vqX3fMMXGynvMh3/cMWZTVPU67bd6mU6Dzpt3ZfdEnY4swIAhyEe39B7xptwzHnr9bR4vKUDmh4tw0MctbFy7egaT/f1fY3l6rhaunt+TYBjJR6hY+YjaU1pFiOKbZ3FY19O9wTA8WreewEAAOiP3o88dvmycPAS60YZn9sX8aOOSNrfEeDt9T4eI7yBcJx2fV37PgDgLZi2BgAgTTwCAJAmHgEASBOPAACkiUcAANLEIwAAaeIRAIA08QgAQJp4BAAgTTwCAJAmHgEASBOPAACkiUcAANLEIwAAaeIRAIA08QgAQJp4BAAgTTwCAJAmHgEASBOPAACkiUcAANLEIwAAaeIRAIA08QgAQJp4BAAgTTwCAJAmHgEASBOPAACkiUcAANLEIwAAaeIRAIA08QgAQJp4BAAgTTwCAJAmHgEASBOPAACkiUcAANLEIwAAaeIRAIA08QgAQJp4BAAgTTwCAJAmHgEASBOPAACkiUcAANLEIwAAaeIRAIC0dDyWUl5zOQAA6IFn47EpTbRtG9PpNAaDwVsuEwAAb6xpmihNidrWiBKzP+u+btOd3I/v4+b2Jn777bdXWEQAALri5OQkBoNBjO/H0ZQmSimP/sw9G4+11hieDGMymZiyBgA4cm3bxv39fbRtG1FmLbjOs/HY1jaGw1k8zuszIqI8N4YJAECvLHdd27YxuZ/M4jEiYn07bh55LKXEdDqNyWQSp6en0bbtbOhSQAIA9FqJ2XT0vPkGzSAmk8nW2z0bj/P57VprXF9fx8XFRdS2Lh4AAIAee8i5tm1jMBgsdlfcZuMBM/O57rvRXdRa4/zTeUzbaZRGPAIA9FqNqFFn4fiwq+K0nS4GCesz89ap8zze39/HaDSK87NzI48AAEegxmxGeTAYxHAwjPF4vNjfcdMuiql4rLXG6G4UzaCJ4XA4C0j7PQIA9N5wMIy2tnF7exsRs+5ra/vs16evMDMajeJ+fB+fPn2KdtoafQQA6LnBYBCnp6cxHo/j/v4+dZt0PI7H47i5vYmzs7MYngz3XkgAAN5fKSVOT04jImYzzE0uC9PxWGuN29vbuLm5ia9fvu63lAAAdMJwOIyz87O4vr6O8f04hsPc4GA6HgeDQbRtG5c/L2M0GsXZ+VnUWqMpTbpUAQB4X7XWaJomTk5O4vb2Nu5Gd4vTM65+3fKfuXT1NYNZJE4mk7i8vIzzs/OIiJi202cvXwMAQHdMp9OobY3hYBhN08TV1dXiTDrZnttpyLBpmogyO3jm7u4uvn//PrsKzWS61xMAAOBt1Fpjcj+Js7OzuPjtIq4urxan5tllIHDn+eamNFFjdtWZ6WQaX79+ddJwAIAeODk5ic+fP8fNzU3cje4iYrdwjNgjHqPMRiCn7TR+/PgR7bSN33//PYbDYTSl2WshAAA4rOX9FQeDQZyenMa///x3XN9cxz///BOTyWSvZnvRkS53o7v48eNHTCaT+Pz5c9SoqWsiAgDwukop0U7b2Um/2za+ff8WNzc3cXV1NTtNz+npXve7dzy2bRslSoxGo/jx40fc39/Hly9f4vT0dDF/DgDA+2nbNk6GJ/H799/jn//7J/773//OPnZysvfZcspff/3vzuOV86NymqaJQTNYHHH97du3OD8/j9FotLjEDQAA7+PL5y9RSomflz/j8vIySpQ4Pz+fzRbfT/Y6bmXvS8XML084mc7my9tpGz9//IzpZBoXFxdxenIa19fX0dZfw6WllNmfKBuvmbjKPpQAwEexyyWg27aNQTOIGjXG43GcnJxE27bx6dOn+P79e1xdXsXN7U3c3tzOzs09mJ12sUaN2PN4573icf6klqOuNCUmk0lcXV/F+H4cn84/xbdv32I0HsXV1dWjeJybH7kNAMDuBoNBjMfjaNt2dvBy08T3b7NTKf79999xfX0dtZ0N4jWDhwObX9heB71IdWlm53y8Gl/Fzc1NjMaj+Pr1a/z5558xHo/j6upqNp1dZ082BrvVNQAAv0yn0yhR4uLiIr58/hKD4SCur6/j58+fcXd3txhtHJ7Mku8Qs7kHjceIWUCenZxF0zRxcz0bJv38+XNcXFzEv/741+xs5teziByPxhERixIWkgAAeX/88Uecnp7G5H4S1zfX8ffffy8OiLn4dBGT6eHPgrPXATMRT0Nvfh6h+ceXPz8/j9D5+Xl8+vQpLi4uYtDMrpXd1jbG4/GihJf/ru3jjwEAHLtFSzXl1/EiD8eMnJycxGAwiGbQRCklrq+v4/b2Nkaj0WxqessR1J0beVwXlBGzk4rXWuP+/j4mk0n8+PEjSpmtgOFgGJ8/f46maRa3Pz8/X3s/AADHbnUAbvkc2re3tzEaj2I6mcZ0Ol0cgDwPzHkzveZs7sGnrZctL/jyiORgMIhaa9zd3cV0Oo2flz+jKc3iiT86Eru+fMdOAIC+mI8yLv//3Hg8jho1ToYnMRgOFh9/i2ice9V4nFuEY5SoURdP8PTkNMrp7HNtbZ89jY+RRwDgo5j30GoIzmdtl0+DuPy5t7J3PG4LutXPPxlRjFkwLg8qikQA4KOrtc5mXbdk0ab9G1+zqV50betdCEMAgP57s3gEAKD/xCMAAGniEQCANPEIAECaeAQAIO3/AcsWUruQqaqaAAAAAElFTkSuQmCC"/>
<image id="image1_349_17" width="645" height="337" preserveAspectRatio="none" xlink:href="data:image/png;base64,iVBORw0KGgoAAAANSUhEUgAAAoUAAAFRCAYAAAACbtdwAAEAAElEQVR4nOz9aXMkSZIlCD459LQLhx8ZEVnVnd1LQzPdH3dp//+PmB2a3aHdqsrKjAi/ANipp4jsB1EWU1U7YBcANYe+IA93GMzU9BBhYWF+/Jj967/+V4MePXr06NGjR48e7xr8rU+gR48ePXr06NGjx9tDXvqAjDEAgDEGxpjG65xzGGOgtYbR9veM29frn+Ws+XOPHi+B+vg8BeeMz3O/+1Booze+r59XPXr06PFyYGDI8gxRFCHPcggp3O/IN9q6Bpi1rSbfiDHW+Axj7EVt+MWdQiEEGGMo8gJFUcD3fQBAURRQSq0vxgAGBkEQbNwgBQX0Se0eL4z34hTWjQmAjb979OjRo8floLWGKhUylkFp5QJgAFxAjDbsu8AMg1Ya2mgwxuBJD9KT68BazaZfEhd1ChljUEpVPwBS2guQQiIchpCeBGMMvu9jEA8QBAHyPAewuUi+1qLZ4/3iuUm5D4wxMJw+Ic/57mMxHo1dNB4AnqZPr/bdPXr06PHeMBlPIKRAWZRgjGGVrOwvzDORQgCe54FxhizNkGUZkjSxQbaycP4VRQtfwk+6qFNojEGe5TDGIIoixMMYo9EIggtobT1erTXKssS3799QFiWUVhvpYvKo+0hGj5fEe4gUAkCapg2ncDqdvtp39+jRo8d7Q5qkCKMQi8UCYRA6p9AY4yKFZkc6tCxLANY5lFJiMBjAu/HAOQdnHLP5DEmSIMsyd8xL4mSnsM4drP89uZlgOBgiiiKUZYnpbIrlcok0SWFgUBRF4zNGm0buvEeP1wJtRk7Bvkn90t/9HLLcGgsyKFEYYTqbQmuNyWSC1XKFUpVuLjLGXvR8evTo0eM5GOyOnnUdnHHkueUODuIBBvEAX758wXw2x93dHbI8w3Q6hSc9aP18logxBrB19pVzjiiMEAQBJpMJfvnlFwDAYrHA3//j75BSggve2PyfipOcQiEEhBBIVgnyPIcf+BgNR5hMJvA8D6vVCv/8/Z+YzWYwxkBwAcq0CSHcTTHGABwQXIALezFGX+eg6HF9oIj0STDn7dDO+u5nEEURhBAIgxCD4QBKK2ilwbjlpVDqQXDhIvX9hqxHjx5vCQZ21kb7LcEYAxccvu8jiiOUqoTRBlxwW2SSH3eserZUSuumpVmK1WqFh4cHBGGA25tbjMYj/I//+T/w7es3PD09oVQluOBnFaOc5BRqbdPAQggMh0OMJ2MMh0MopfDHn39gOp2iKApwziHE2iEEYEOgtaigq7ShC+gDFj0ORHvQH+qkXcQBYjiLU/iSEFxASIEwChEEAebzOZRW8KUP3/fBOIMwAkbUqtle0Ent0aNHj2dxnf4gALvJl0IiDEMM4gFWyQpKKwghLEewUl8RUoDpTVu7a+0yxkBKCQbminWFFFitVlgul4h+RPjw4QOGoyGGwyG+fP3ieIda65Ocw6OdQmNsClgrjcnNBLe3tyjLEv/59//EYrFwqWBPerbyURu7gPL1ydVJki9FluzxftAY9AaNTch7HFulKsG4TTvkWQ5VWiMhhXQReQLtKnv06NHjObRt7UUjewxX7RgKaR1Az/NQzi0vkLKqgN2sn4JG8a5nXTZSbSnLEv/8/Z+Iogj3d/f4l3/5FyzmC6wS6zSeUqHMDu1oUi+DDoIAcRxjOBxiOp3i4eGh8b6tX1Q7sX2VM+9xEe9xPNrjCbBRaAYb9aqP10M4HD8D2pO/fl/GozEGwwGMMfjy5xcYY6C0amzOCP0c7NGjRx1t2+I4yKxpL4x+XmrlZ0I941mPyvm+76KGXHB8//YdeZ6DMeZkwk7FNqUWrTUYGKI4wl/+8hcEQYA///gTi+Wi4ZgegoMihfUUb+AHuL29hRAC3799x3K5POJymsfr0eMSIHkYmpT0h3MOow0UUw0JgPc2/jjnALNVbapUjfnMGYfG+zHiPXr0OB1ka8mm1O2tMQZaWXWR9+QYboMQAjBWn5kp1tRovjBorQOA1XKF/9//9/+HX375BX/55S/49u0bVsuVTTvzJpVvF551CskL5ZwjDEOMR2MwzvD121dMp1MIIS5S8UK4FpmPHm+PNh1hG8ePcQbJJVSpoIxqfO69IEkSGG2wFEtkWQYp7LTvK4579OhxLKgyFthcc7nglq+sTqskvtb1v51WT1YJEiQAgyvk25aVcR+5kDwaFxxlWeIf//gHjDEYj8cwxiBZJc6Pe84xPMgpVErB8zyMRiPrEH79ivl8vpXE+JYcwZ6f+D6wjYoAAxhmbAXbjnRou7jpvcDzPMslNNjg7FxrtV+PHj3eCJVp1Vpv2BMhrZII1zYDcYyt/Vk26/UgGXUu4eDrimLTrLK+5HpEzUFUaYt+b29vMRwOwRjDcrG05/JMMGCvU0hRQs/zbISQMfz48QNpmsLzvL0ndsrvzsVL9wTs0T1QpNqlRU21OYBxk5OE04Gf2yHcxSlkYOtik6rLELDbIeznUI8ePbbB6ZpyDqXUhj31uAdjjKPuvCYumbE8FRuBKQZw8HWBn4Gj65y6Fu2zz3UOPWcc89kcQljtRMA2MqCq5F3YexeNMRBCYDKZYDAY4OnpCYvF4pTr6NHjxUBOIPk4xpiNVPK+tkI/K8hJpk5C2tg/pvqv30T9PKhYtW99Gj3eCdq2g6JP752SQpFBbTSUVlCq9Ucr19HkRcHsH6UUvnz5giRNcHd7hyiK3HnuwtZIofuAAeJBjNFwhK/fvjqv8yW5Av0i1eMUUFUXFZwcsj6+JX/ltcY559zKGLSkegjUdvK9Ocw/E+p82v459nhpvHS279rBGIPv+Y3XuOCO2qSUQlEWLzZXG/eQA9xwfP/+HYILjIYjZGmGUpU7P7/dKdQ2kuD7PgbxAPP5HNPp1BqeA6/jZ3i4PboPCpU3ZGdqVXEULbs0usxfZbAO8nA4BGccURSto6kAYGC7nGiNLMtQFMXbnnCPk9GOEDp+bc8V7fFCIKkvx9XGukPSe4aU0vUrDsOw+TshbX5GG6xWKxSL17G51BFFK43Hx0cIKRAPYiyXS0spYpu+2s5IoTEG49EYAPDt+zdnaFxpNWuGkDeqP+vf0xupHi8A2nWRuCdnm5VVLxmq7/LGhzOO29tbq6a/JURYliUMDPL8iP5LPTqFts11G6HXSE/1eJcgweQ6qKLVkx4MTIPD/V5gjLHFuMMRojhq6AIyxpzig4FBURaOk1l/zyXPpQ3GbUeU+WyO+w/30FpjPp9vTfdvLzRhQBiGCMIAX79+dST1bai3rasbKOJ40d/a6N457PGiIK4cx7pLx3szUAzr1PlyudxK9+CMIwgCBEFwlKhpj26A7OyGs0+7/ivvDNHj+lDnddOm5D1tTLTWyPPctbejfsUEwQX8wEcYhPDk7iLdl0BddSNNU6RJiiiKkKZpwzElbHUKGRju7+6RpZnVIqyHhSsCI4EzDs/zmuT+msq5Vtpxvdrq5z16XBwVd46BWVLvOzNOgJ2T2mhMn6a2d6YnNyR67u/uEcfxuyeGXyXYOmXXeHlLG9EePV4TtN6/Jxhj08J5nrs2wG0ON+cco9EIvue/eJ/5bVFHeq0oC8xmM3z+y2eMRiM8PT01JNsYY9udwngQIx7E+PL1S3PHyWq7VDJA3HZFUEY5XhdVNkohN1IZxHnZhT6S2ONQtBc+zjl833cciqIs7IbkHS2QBpUuViXPILjYaPNH96Ioi4MKcnp0A/sihO2fGVhvS3tcHG1bKoSAlBJCWDtDMjWvLVz91qjL4WilN6P1lUYs4+yo2oxLgp5dmqZIkgSj4Qjz+dy136P7v+EUMsYwGo6wXC6dHqHWeishsRF90AalKm0VaKWcLaVcRxarm1BPb23De1m8e1wG9TEohIDv++CcIy3ShjN0zQbnWND8C4IAvu9vFNswxuD5Hoq82Jo+6NFRsC0OIZ63qT16XBJtKRopbSai3t7uPdlbxhi4tLqMvu9jMp5sREs5sx3hGGPI8/zFoqnP9bLnjMMYg8VigSiKEPgB0iRt0IgaTiGJTnqeh2/fvm10gtjWSYK4BG7haW9iK65hv2vt8dIgErQx61D+ewRdtyc9hGG4UWyijUYQBEiSpK88vlLUuYMGm7qcPXq8BpRSUKVyTuF7hRACWZlBCIHxeLyRImaoqoArCbA3Q3VaeZZjuVzCD6rMGjnzqNLH5FlS+XKe55jPrSahUmqro1eHMabh9O3qQ9ujx0tCKWWraY2trmX8/YozG2OQFzmQAGVRNuawFBKlKKGU2kgt97gO1DncRhsbRXxhrlKPHm1ooxsZQuB9RQmBtQoG57bv8HQ6bXZ8Y7C0Jk9CaYUsz97uZGGfT6lKrJYrTG4m8HwPWWbPycCsI4XkFI7HY6tho7Zr2LTf7xYV8glNkwRNCt8uffzOBkyP14MxxlXKv+eNCefcaRASXwRY35MgDGz6uHg5AdUel0f7WdV/NsaAM6sE4TbpFEXsbW6PF4Tj0OF9ru+MsYZT+PD44CRoAGuP40GMMAxRFMWLy4C1U8fbnolS1jk1xiCOYhs4qN4v6x8WQiAIAjw8PIBxBq30umdf+4ur/4w2m/nxujPp9HLXQpc9erwU3Dh751GTeg9MAlUaRywCA+udwisEje9tz43Xupa2szc9erwE6lI079EhJBCXTyvbRlSrddSU+kAbY5Bn+av2hN5ZZFlJBymlXEW0UgoMzFoR8nR9z4dWGmmaQgoJxpm7gDqHcFv6mN7j3vuOU3c9erwlnnP0gjCA0qrnE14ptorT9ra2xxujH4Pb1VMYY/AD2/YuSZM3zWJRZTgVluRZ7s6HCoo5YGUriqKAkJZDWJYluOAQXEBp5Q7WOPAzu9BGL85+w9qjR2cQBqEjPPecwuvFtkX4Pepy9ugGtmln9rDzNPADAECapG8fwTe2MAbMcu/rfOSGTqHWGr7vO6HpoljLVVBeuhERbHUnoQo4xhk86UFIgSzLesmLHq+Ctjj6IcbpZ108t0lHaa0hPIHhYAilFVarlavU7nFdaKtAAC1aTv9Ie7wiVKkQhIHtqf5O1/sNm8utzQ2CAOPxGFEUYblcIi9yaK23Zlxf+twoQEeFMXVdSd/3UeSFTXcDa10zKSRUqRrSHsRD2hYprP9XPwHG1/l1bfTbe8Y9fnrQpoSaknPGHe9113/vBVprSCkRxzGGwyGyLEOaWh3HPlJ4/XALTK3FWI8erwUubNMAxnvpOUJZlpBSYjQcYTweoygKLJaLN7W3TsYKcM6g1hpGG0sXrJxHTm+QQkJIgVKVLmVcV+k+FFJKV4Xz3trd9Hh7eJ6HIAhOGrs/K3zfx3A4tG3tOHdVyT2uG4yx9eanFg3oncIerwnf93ub24LgAqPhCKPRCJ70sFwtsVwuwRl/037zdcfQ2QnW3FiuI4ViHSkE7EWdEk2htlp9ZWOPt4CU0nU16WExGo4wGo4gpUSSJlZRv48Q/lSoO4N9tKbHa4ExBs/zdtrc99pbfTgcWoew0gCcz+dOL7YraxO1RK0rxDidQpKd4ZyjVCUEX3uyG8rcOzRwKKW8SlYA8G6FLHu8Hmj8CSEghIDRtiMPkWi11k6n7b0aJ8D2MjfGIFkmSLPUaRfu0rDqcR2oF/y1aT79hrzHS4Ha2hVF4TbhMPZ1KWWjBsFoS0F7T1lDxhh+++03lGWJxWKBNLG9hrXR4Jpvjea/ph1mjMGwLQXAVUc66xRy7iKE9ZOtO4S7iJHthaWPQPR4LXDGbYRbSkhhjZEUEpxx+J7vJp9W+l0vkov5AmVZIi/yPm38k+I9Lbo93haCC0hPug5oQghwYdvjEk9Za2tzc/X+7I0xBk9PTyiKAmmW2qyptpx3bdb35s035GY73UTuePtBDmGPHm+JIAwQRzGkZw2T4AJCCisBEAQoVYmyLFHkBfIit3IA79A5nM6ma1Jx1d+8n9M/D9oZmx49Xgq+72MwGCCKImijkaUZPM+DJz1opRGGIVSpkBe53Yi+w00oZxzfvn0DACitXEvKtu7zW6CuIuNoJiRJw1odTdow2jQcw054tj161EDcODJKlDYG1pMuz3OslitkWebSHu8J9Z0g5/zdpXLeC3pnsMdrYLVa2Qp3VJtLzmyRqrAbcnIEkyR5lw4hYKP2jdqMjhaB0fkcFCl0b9LYcAyB3V5u/QsoEtH+Qo3trbd69DgE9UpLziw/I8syZFnmyv9LVeLhx4Nr8g2g2aD8HaE9V3uH8OfDe9vo9Hg7eJ4HpRSmT1MAgPQkojCCEAKL+QLzxbxTjs9bgebkPnvbtXlLgb+tTqE22kod8GZK4rmLoEgEHaPnF/a4NAxMc9MC21uSdq2Nvts9evTo0ePF4Pu2fVvfHekw7OxF3CFsDdNxxk9aWI0x8HwPURTBk967Egju8fooVQlV2ibenvSapf4M6Idfj/cAqq7vsy49XhtRFIExhizPGvImPXaj63zurVbknBOWUsLzvQZxsUePlwAVTwBrmYS+o8MmGs5Cf2t+avQb8R4vifr4opa22qzbpfUamdePvVvLNj9w7/uqsUDl18YYpx/Xo8dLgFLGXHBEUYQiL7BcLm30kL2vVna7QFF/zqzsVFmWb31KPS6EekcT+rlNau83SD0uCc/zrAas0bi9vYWBgSoV4jhGFEadjoC9Bihi7yL35vrm4s7qY+B5Z5AWXup37HSLpLCRGzAYblCURc836HFxCC7g+z7iOIaQopEu7h1CC+oJzRhz/B9qY9mjR48ex0BpBc45wjCE7/nIi9wqGiiNoize+vTeHFRYQpvx8WQMVSosV8s3PrPDsTtSeOCayjiDkFYjjjNuteK4sOR/wZ2DyDnvF+oeFwUXHGEUIgptlLAoakapH2oA1tF+uldBELzxGfW4NGjzTpSdxmvvPHLT47LQSkMIgUE8AADkWe42mXmeX0007DVgYHB/d4/JzeStT+Uo7BavPsCgGGPg+z6Gw6H7TBiGCPwAnu+hLEukaepSy1rpPkrR42wwrKuMObOtGZerJYqiQBiE7n3aNDuZvMeUMmPMaYpxzgFu0+7XlM7ocSCcFi3ruV09Lg7yB0gTNk1TpFkKLmwA6L0POdKANca4DVocx65ZAAAnZN3l+bk3fXwIyrJElmUQoooIMo6ytFWhaZqiLEuXwqKF/L0tzD0uhzpdAQaYL+ZuAyOEcBXI2+gK740IzZmN1FP7PwBQpUIYhiiKws5NY46qWn1v9/Aa0Nj4oC/w63F51KliWZYhL6wwNcnQCW7X/zzP36V9IBtKzl8YhbZ7STUXw9D+XKoSMOtOJ13E+U5hUWKplvB8D2EYolQlOOeuzyotPK69S+8Q9jgTBgbQgIItKKEhNR6N4fuW50L9jtuRwvcCzjmEEPCkhyAInD4W5xxKKSfmTZs2Qj8/fw7Un+N7XKR7XBgGMMwWlCqlrEYsYxgMBgjCAFmWvesNI7WwC4MQg+EAo+EISls7q0ONu9s7KKWglMJ8PofKu5sxPdspNMZAaQVpqhZixrbI09qWqWul3ft69DgXBtYwOeNTG1ZFUbg08nsubOLMpoqp6IsqBAG4gjDOuXMM61xMg+Mihz26g10boN729jgXZHfbHTqyLANjDGVROtvyHscb5zZ1HEURPn/+DCkkSlWiyAsYY3B7e2tle2CwWq06nUI+2ymkfDln3BWUGFinkKRp+khEj0ujbXgYY1iulmuaQvVfVyfeS4MihZxzpGkKpZR1FgV3TiHN2zb6+XoloOhNBXpW73XM93gd1G3varlCWZRQSrkitvcYpaZMKOccg8EA3759s/2fq0Icz/MwGo0wHAytUsZbnWfVyg7YnTk72ymkg3ueBymk20k4sqVe37B9J9KjxzHYtiOlDUh9cXyP441EvbXW8D0fqlT2Z2igtNHCIAhclH/b5+t4j/fwGkDRG0KdzN6jx0uhbg8YZyjL0nENaVNOeC9jUWm76SauZZ7neHh4AIO9P37gYzAYoCgLxzV8LX952zPYVdvBGNsvXn3QF8JASIEwCsEYc2mqHj1eC73T0oQ22lb6V2LV+wzzezHa7wHvmdPV43XhJI/6TAKAyo4ecSu6vGad7xQagyAIEAYhsjxDURa9PlaPHm8MonCUarODSXtu1hX3eyfxemHQP78eL4t+XT8O17hJOzt9LKVEEAQoygJpmsLzPDAwV+VIujw9elwaVCwhpR3G9c1IPYWcrJL3p49prCzPtsh9I814fTarR48ebwSnalDZXdcKt9Zq0RiDxWJh7bFpbUB/YoNjtEGe5/jy5QuWy+XGJjuKIpRliTzPO10IebZT6Ps+OOdYLm3Vp5TSPXitNWD63UWPl0EYhhiPxwiD0MmtML4ea6pUUFrZftz5Jn/uZx2XJFittba9jhlc8Q3tz+h3XTZOPXr06BYYGIaDISaTCaQnN2wIZ7bQNMsyKK02ncKfOJJtjEGe5fjnP/7ZLNarWoyGQYhv82/I8qzTvO2z08dlUWK1XCHPcnie5yqQtNINJe8ePS6NespTG72ueK/+cGEr4kma5T2ORacRSt0uKpFvrS3vsC0x0aNHjx67oI1tcyc9aaXnVNPmGtguZ0EY/NQO4DbUg2F0P2BsdHU8HiMvcqyWKyfT11VcpKOJUgraaIzDMQLfDoaytFym96pb1OPlkSQJyrJ0avGMMdtuqcLt7S2kkE5tv9Eb+R1gm1adS6tXFco9evTocSiMMZgv5sjybJ0JrGVnJpMJBoOBFW1W+l1uxNsQQlinMM+RJIl1rPF2sjTP4Syn0HGTKg85SzNM9dSGUYu85xP2eFkYG6lOka75hMXaAbq9vQVjDNqsuXXv3Ugxxpyo/M/M7+nRo8floZRClmauQYDrqV5hPB478fy2ZNJ7AK09XHAwWFt7c3MDz/MwnU6hjYYnvU7b3svoFFaFJWVZbkRjunzxPa4bXHBIIeF5nuvxu43fYoyxrZl6OKOlte4j+D169DgKRhtwjyMMQ+cU1iH42g5zzt9dNoL8HaUUPOnh48ePuL29xXQ6xXw+d+nkLhc+nuwU9hpFPd4aQggMh0O7O63aDNUhPemcn35zskYvPdOjR49TEAQBhsMhBsOBixLWsy+cc5SqRFmW8KSHLM/e8GzfDlprZHmG8cSuTT++/0CapShV94v7LpI+PhSO1/TOU3g9LgOqfJPS9t3mpll93FDe7zcwANaFJ32BSY8ePY6FUlbRgTFmC/hEs4CPM5sxLIsSUsp36xQSh/3h4QFBELhWo06mr8NazqdHClFdVNWuhRw+xyNgtfegqbZf5xp29cb06D6MMVgsF661EBWUGGMQD2Lc3t4iSRLHJ6R0cv3zPzO00RtzELrZ/7JHjx49DgYD0iRFWZbgjDtVh7IsMRgM8OnjJ6hMoSgLt1k/GObnoZspZfsdz2YzDOJBwyEEuu33nB4pZFXPY9+zxMnqYqWUlmRZXXSWZcgyS0ytL0b08PsITnfR9cpxKppIkgSAdXaklOCcIwgDaK1thXKtq8d7a9Ze7wUNwMn39OjRo1uoC+53FYwxaK2RZ7n7WUiBsigRRzEYY26tL8vyqPXdsJ+rMIVzDqMNVqsVlLYKLV2OEBLOKzRhVqV7Mp64l9ocgyzL8PT0hDzPO38zejyPuuHqmhEjXSghhO2yUxQubC94dyUAevTo0QOAy7w1X6rZ3I5t1IuiANi6uxRtxBljyPMcnJ0thXyVEFzA93xEcYTFfAGtr8MhBM4VrzY2TFqWpSWXVgRT+qOUQhAELqV3DTekhwXDnkIi1vq7I6Cm5J70EAYhiqJAWZZ9oUmPHj26D7Yjc8baP3bH8JK8FePMdTNL09TK0uX5W5/em8HAIAxD/Pbrb7i7v7sahxA4MlLYuKgq/79arpCsEvd72i1wznF3dwc/sG3wwiC0jqLpbil2jzXfk3ErM+RLv2GUtLLVvEIKqFI5kfK3hjEGQtjd2XA0BGOswSd8zzgnXUySPj169HgZuMID2G5DvmjaXFUqJ8xfFra4bp9j+Jr0EC44uOAYDocIoxCLxQJaaZudEaJxLnV+83vAaDSC51t9Qs65bcXKbDFklyXBzksfm9oArDiGKrXVSVEYOe+Y8arTRDf8hx6HgK2V6hmYe86UwuCMQ7NucNOcYCjnCIIAcWy5LdR/k3P+U3FVevTo8fPBFW5WflO9eJMzbh2KjjlVjDEEQYDJeILAD/D09ISiLKCU2tAwbPObf2ZIKeH5HhhjCMPQ+UJaaxRF0Wnd3JOdQlcoQo5DddFCCEQyQhiGEEI0+tP2Kbzrg4FpVE0BdnfYSCF34LFKKRHHMSY3E4RBiKfpE9I0XQusduAce/To0eM5OG1Vsrkdtl1xHGM0GmE4HGK5XCJZJa7QRAr5bovafM9HGISQQuLzp88oigKe5yFJEjw8PjhaUxdxulNoDJRWuJ3c4uPHj+41mHXVqjbacQ61tv/u2k6nx3ZQqN8Y0+hSwzm32lRgnUgt0vdHUYTPnz5jOBxitVrh4eFhTXTu5tzr0aNHjw0YbTfiVK3aLtZo2923LOb4+OEjxuMxyrLEly9fUJSFK6p4rw4hYIMUvu9DCIGb2xtoreH7AebzGVarFRbzRWeDZEc5hW2NHWpnUw+FMsbcIsxgw6VaValHbQC+/vx7rUy6KphNXTvGKodQv+2gpirjOI4xHAzh+z5msxl+/PiBLMv68dWjR4/Ooy3TVocxBoYZMM7cH7Qyj6/pfHnSg+d7kFLi9ubWacF++/YNs9kMQq5VHt5LcWndLzLGQCuN8WQM6Uk8Pj2iLEssF0tMJhPEgxhhFG59jl3B2b2Pl8tlo9hASgnObHn63f0d0jTtdKi0xzNgu4U2acf6VhM/yzKUZYkwDOH7PpI0wcOPBywWiz462KNHj6uC0QYatpKXaDm7qlbr6+lr2t80S1EUBUbjEaQn8ePhBxbzBWaz2btwALeBrpuoSvHAptSTJMEff/zh/J/haGil0czPKl5dgTxjQlLYSuTRaGTL0rMcRVm46ilCH8XpMPaMV86qfpcdIAz7vg8GhtVyha/6K8qiRJIkrpNHjx49elwLTPUfM6yzm9oojFCUBebz+VqOrrBydBQl7HoAaJ/WY502dUx6V0qJNEnhSQ+TyQSj0Qjfv33H09MTPM8DYO8LSff91E4haRIShBAIw9D2/ssL5Hm+rqJ6J+HknwEuCrjDueoCn5AKYDjnWC6qiPUura8ePXr06DiMNhuqDnVHBXhbpyvNrAah53mYz+bwfM+dI3EJuwzS393p8J1YQOkKbaXAIB7YgFiRu9ar9J48y5EkyZuvnftwtlPYhlIKDAy+70MpZRti13sjV44h8SD6iGG34Ca1sZqEdb4K51aTqi5F9JZGgCKWxGntukHq0aNHj30wqFq9VZtb0rUDsMHffwuQ86OUAhd8fT6s2zqEdf1dIQQ87q2DWdscQFf4fZjzprUGFxyDeIBPnz/hx/cf+PHjhyvU9D0fcRQDDJ3WKARewCk02ip5D+IBlsulFQ9mcCnmrg6aHmu4tkrVRCJtQsEFOOfQRluexBsXmvTo0aPHT4tKK1YIm5bVWnfaobiKtb3SgeScw/f9RsaLZIC01ken710rVWa57rP5zDbrqHRyozgC5xyL5QKqVJ1eOy/uFA6GA4zHY4ABq2RlNYv02xYk9DgO7efEGXcGijNum3sr3dmS+h49evS4VpDIM2d8vRGvVDy66hBeC+rRTOINtot2SF3jGHBuo6bfv33Hcrl0xwcAIQWGwyEYZ1gsFla2p8NyPRdzChmzvQ/v7+8RRiFms5kl/ZMQ5ztSM/+ZQJw9Lqyaftcdwn6c9ejR45pBDiHnVerYVFxD002nkDp1dD7oU2/XWnUWodfrrV2PBUUXBRcQ3DbsSNPU1VZwxhHHsX09Sd+cAvAcLkLo49xe9F/+8heMx2MURWG7SVTOA6Ufe1wf6LlRb07HJ+yebQKw3v0BV5LO6NGjR49tqMyX1hpKq046hCTDopTqdH0ArV91iR9tLGee0vL0PqC5jhxy7DpUqVDk1uEUQmAwHGA4GGKxWCDLs4ZaSxdxdqSQc47BYIAPHz5gMBggTVNMn6ZYLpfI8qyTA7nH4aCJYbSBgnKTqIuRQgPLZy2KAkVRQHDRO4Y9evS4WmitbZSwo1xCxhgCP3DRwg4uCw0Qb3BbNsk5jSdkmtoO8WA4AACEQYjJeIKiKGzquOh26hi4QKRQKQUYe1NWqxWenp6sR1wJC3dxIPc4HPWuNSQ/1NVnGgQB7u7uMBwOIaXsHcIePXpcHerRq7IoXeu4LtrdKIrw8eNHjEfjTp5fHZS13Heel6IeUWe38WSM29tbZFnmGn10/T5dRLw6SRM8PNgmz1me2b6N18Ax6PEs6n2sje4YFcDAtoCC5YIEQYDxeAyllG3MXtoQvjGm06mNHj169KhDGw0ouKxMF2wuRdHqjlUQBJjcTKCUwnQ2XcuD7dMCfEsQP7OlBck5hxBi3cL1zHMvyxLjsXUItdGYzWZWs7nDVceEs5xCxmy5PA0IhrUSuKvi6bhX3OMIdEwYWhsNZhiEJyCFhBTSjr8q3QJs9hXt0vn36NGjxy5oo618CuPdWEdrm3DSTmSMwZNWwJpEmsn2ds0nJN+EOJp1vryUEr7v74zKHuuUj0Yj/PKXX+B5Hh4fH/E0fUKWXQed7uKSNG10YYfT4zLo2rM0xkB6EnEUu046JJw+Go1sS6GyRFEUKMvSOoTduoQePXr0aKAdTOmKI2FgUBYlwiBEHMdgzNrasizhBz4G8QBaa2R5ZgtNq2xhl9YNJw5eA7Xgde3tLnC/byY3uL+/x8PDA758+YI0Ta+mycKLO4U9erwUhBAYDUe4u7sD4wxSWB5hGIYuFbBYLDBfzF2nnR49evS4NtSrYt/6PAbDAT5++OgkXDzP9vuV0mZq5rM5jDZYrVYuotgVtKuKGbPXQNFY0lQ+F2mWYr6Y49v3byiKovMyNHVczCmsC0FuE4PscZ2odzTxPR8AkOe5+/1b8kaEEAijEFEUIUkSLLPlukUUYxjGQ1v1tVw4Adge7xfXuinoJDerx4uDHC4Ajqf/1k6hlBJBECAexMjzHEVRYD6fu9Z3cRRD3AosFgtIT27Y3PZYfus5KYSA53m2ZZ9WUFpdJO09fZoiyzIsFgv3DK8FZzmFNECfa9bddzO5blCpfhiGALAW/QQsz+SNFi3agBRFgcenR8znc9eAXHrWeJHgK2lp9Xi/uGYb9NbOQI/XB2MMURSBgSFJEhSmeP5DLwzaXJdlifl8jtls1iie+OWXXzAYDqxu4TM297XpPO35T61bSalClepicmt5kSMvbPAky7Kzj/eauGhHk10Pud/p9ngNKKUagulb2xf1i2uPHj2uDWy9Oe+SDcvzHKq80s22AZRWyPPcRTr7bNKFnMJ6P0HGWKNKVRsN6N4xvDbsbBfXoWCLMTXSsIFLHe96b5eMaY8ePXociq4UyW21oR04r5PA1ml5p5xygTXi2teZs51CrTU0tNOJu7u9g9IKT09PKIqiu3pFPXbCGAOwddpfSMu7kJ4lEvu+v269pDeruV7zPMuyRJ7nKFUJxplLbfi+D8aYVZDvG8m/GmjMcM5dH1ESP+f8NGkNt+GsLYxvnQquf7+7Jrq0badmWu/t0QNbUppVgIVsrhACMICQYt3dxLxhRyljHanVaoUss5rEJEsnhXRdzbS5Ap3iivrUziidf1jj7GDXIruH4GynkC6cc47AD3Bzc4MszzCfzVGy7qt399iEgYEnrBMopf0jhIAQApxz+L4PVSqUqnTG4U3O0xgsV0sUZYEszRoTms4xz6zD2ON1QEaQUvk0fqSUEFwgiqPjjodaBqL2HadEJy5li0injZxdVVrNM6Vtz9NSlVvTUPWMSm8XewBwmwXGrVYeOYI0Z6gy1vM9W9iRF0iS5M1smjYaWZrhUT+6DleCW8fVD3x4nofv379fRfOKl3KsOeMAX2eyqHFC19vbEU52CttGmgx1URR2B6HVemf/hsUIPY6HMQZcWOfP93076el3VVcT6nDylo/VGIMkSZAkie1qIjgYGDzPQxRFtgdyJUYKvH106T2BMw4wIIojxHGMKIogpUQUHucUtnFO0dolHTEpJQyMSz9pre2CnSbIsxxpmrrxV//u3hnsUUddVN9VwnLuNhBSSjuXFOBJz9rcNzRjxhikWYoss5twzriNCnKG4XCIPM+xWC6glQYX77eLFIPlKJJ+42q1QlEWVzH/z44U+r6POIrBOcdgMEAURzDGYDCwDaGp31/vE14PXNpVa2RZ5nawnufZFnJJgrIsbZTkDSt6ySgxxuwuzNgdtyc9hEGI1WoFVaq++v0VoZWG53mIBzHCMMTd7Z3l7pS2d/bT09PRx6w7VCQ+e8om85IGuSxtpMbzPPi+j7vbO4xGI2hlaRVlUWK5XGKxXLiNclmW10vK7/EicHbJAGVRuhQxGBDHMTzpIcsz51SQ3X0L0Pwh9QkpbAaJ1B2Gw6Gtks6vw/m5KKrgFyFJExhtMLmZ4NPnT/j+/TsW88VVOIZHOYX1YhKKAoZhiI8fPyIIAlvazRmGoyGCMADnHMvF0il699HC6wFFQIqiQBiGGI1GkFJiuVxClco5hG/pcDUKnKqddlmW8HwPRVEgzVKUquydwleAMcaljIajIf7yl7+AM+6U/N0motIBO9oWbOH/HHNu+35+7nvbnzUwrrG9lBJRFOH+7t5yXFUJIQQGwwHCKMTkZgKtNVarFabTKWbTmeu0Ux+7/fh8p6gVx5WqBFP2B6LrSCldxDnP8ze1uUQNqVMgKI39+fNnxFGMr9++ug3TVaSQa7J654CBuawURXhh7PHDMMQgHmA2nTknusvyaOf1PobtIuF5HpRWWEwX0NpGChhjCILAdZcAer3Ca0J9A0AGioGtxaG7UHLGmgu80gqDwQC3N7colS1A6WKrpZ8RnHFwwTEaj/DX3/4KKSUenx6RZ1arq2F8W7vqg1CNuYs4hcc0pWfbnUgy7nXqDBU5Aev0OfWDlUJiOBziw4cPmE1nmM1nyNIMaZba99dShj3eDwwMmGkqdjDGID3LJzQwTox/G7/2LVDvJ+9JS9UZj8coVYkkSVyRSdflXepFcfTzqVG8UpWQUiIvLIc9kIHzfwI/sM+w6gBDNqKruEihCWDTxD9+/AAM4PkeOOO4ub1xDuI1RAmJEHpqROJnhBACQRDY6CBTnb4vgR/g/v4eQgp8+/7NGqgr2K1eM4wx4IzbiFkc4ddff4WUEg+PD3uN3yHPpMtjbQNmvaiQoHodQRhAa404inEzucF8McfDwwMeHh6QJImLQDL6rx+z7xaMMdcFoyiKRlV7vcNUFyClxN3tnd0EPj46mwus50NXzrUNBhvRC3zb5CBJktOPVW0MgyBAFEXI8xzD4RBhGLrnFQQBAPz8TiGBokilKqFSKz9BnC9ClwdIHe9dRqdeRk/kZ0oTNO5Lx24R4zaEP1/MXdqyjxK+AhggPWn7nwobISRZoDzLT3burlHOgdBuSVYUBTjjlmtkDG5ublzLsB8/fqw5h0o1JS26EJHv8apgzPKiAThZN5gzouwvBBdlY8BiscDj46OrH+h6cZ+TWxMCfmAl1s51CrXWuLu7w19/+yvyIscgHsAYgyiK8csvv2A0HMEYg6/fvuL79+8XvJrL4iSnsO7cMW7lGbIsQ5ZlMDAuFcIZR17kO0ux6w7jW6J9HmSMt/Vx/tlBE51oAKPhCL7vYz6f2zZ3BliZVSfL64uiwMPDwwah/1K8kR6b4IxDCOEqjOfzuUsZ53m+ce85jpNnaOsB7nuGuxzItgwM49XPz6SRtx3P2Qa2vq5tdqwezbELRgnDOGhFT9MVfF/i8+ePGI2G+PPPP/Dw8ABjVO0aGcBYZ5yAHi8Dxi0NqygLMMYwGA4QhAGyLHM6hQBcNHrj863Nw0va5vb8y/McX758cfxzoBlU6coa30ZdSo98Fd/3XaGYMeaoiL02Gr7vOw6oJz1kWQY/8EGHIK3Jrq9DFxGvLorC8guq6lSgSiELjmSZdJpUuQvvNVpI2kqe52E0GmEwtGKkRts0oULN2erQ/dFGQ2XKLcZdn3g/C7jg8DwP49EYRptGauQo7t4B6FLk0KXxdkTyGkVQnMI76+g7sBb1DsMA//qv/4rBYGCrFBeLzlxnj5cHFR540lbtR1Fk6TqlFYZ2toxtnwNvGU2mOU/FFcYYK0fTUWcQaAY+6pqnrpLa8JPWNlUqTJ+mWCwWkEIijELc399DCokvX75gNp/BGIP5fH7hK7osTnYKiQOzmC+QZZmtkCoKm26UHuI4hhACeZY7WRD63K7d9VujvrNvRzjem5F2GlRV5SRgnUDaRXUNnHEwbx0B6mIk82fFcDDEYDDAbD47eAN4yPy/Nm4vZRaobdZzqNub0Wjk+NcArJySu5enLfrXJpr7XmGMgTLKdjGRHmCANLXKCTbS1NIE7gjnlNZJrXQjXdzFtZ3AGIPv+wiCAJ7nIfADeL4HY4zlzleqGskqOaopA2fcSlFlJfRKI4ojjMYjxFEMz/cdZ5GKWrqM053CapdcqhI6Xbe5I82iKIwguGg4EdfCKazb4LqDeDXnfwbqIuSLhXX40zRFGIZgYGuuVMfWasYYbm9uIYTAfDHHcrF0UcP38NzeEje3NzZS+440+MhhbbccM9rY1HJ9uGkAtXSz1tq1/OOcQymF5XIJALi/v4fv+/jzzz8xn88bjuGh47jLi3KPTdSLk1bJClJKZHnNIXGBwm7ZMGMMfvn1Fxf9Wi6XnTvHOkgtJYoi+J6PsiytbmDlyxhdObhKu3l9yPXQpktwYSuMA1tPIYWNnCarlX2+eWEbLHR8LTrKKdwWPTNmXTKvtQ0be54HP/CtU5Fm6xx9La1HN/KtDRhVBGVZBsEq6RxtO3oIJmyUs270f3KOoTHGRdqSNEGSJggC275QCIFVsnJdTYC3uQfbdsqMM0RxBMYYVskKQRA0upkAm2Otj6CcjzAMIbiwFbQwjq+3E0fc8jaFg2zNxbDP9BwjZVg7L2NsNJ0WhPWmpGk76uOSMeacP8YYxuMxfN/HP/7xD8xmMyiloWupeM645XJvoUnQ/K1/1zk29tqitdcIeoZKKZt6lBJhGDqe7mq5spvxalDWu6C8JUib+MOHD7aLWamQZRm00Tuj1G+53lMHoul0CsBWTo/HY3jSwypZuU0YaUHSZ4BN3mYdggv3ftIvHQ6G+OWXX5Bmqc24VVzF+jG7istUH9cMooZGPIgRBAGWi6W7SUD3nShyEIH1AGKcgWh07yXi1J7IxhikaQrGGIq8sLuoN1wo3EJVaSaSJApN6LIsoY3tu0u8LQANY9XjCtGhykuYdVSwHjnXRoMbvt70kudZs4HPiWmT4O2vv/4KzjmenqZg5BBQdLLcXnAAvP1Gu8dpqAdblFJWgD9Jrd6q0a6dImf8zR1CwDqlYRBCK42yKJFmqQsUlXrdNKBLKVOal8SB5NymfesZsFOkdFxLP235+MPREIwxTJ+muP9wb4NMXIAL7igmXcVFdAqpLB2wrXk+fvgIAFgsF7b6uOPl6btAO/FrO+9LgjEGrTTm87lTbe+Kk08yOb7vw5OeS8kFQYDAD2zDdlVaUrF6W0f2Z0V9jmwbD+/lnjNuAKMB0DhbFwe0/tEA2cb6wkmcxOFwiM+fP8MYYLlYV/zX6Szb0C7weS/P4GeBK940BlmaudZ3ziHs0HoURqHV3xzElpunbQBhlaxQ5AU833vrU9wKzm21sed569aCJ8IYA8GFez63t7f4+OEjHp8esUpWuClvbJtPVUIY8fNHCus7Fs/z8OnTJwRhgN9//x2LxeKqHMI6sZRx5sLC79moUmPvoqzkBrakq97q2dafjZACYRACDK6pPO20kyRByUpnaHv0OBXbHDKbGm6OR2M0WFWoRZsVYN36i/iE9DppapJzqI11DEajEbQ2+FN/QZ7ngLFVkvuiL6vVakMnsUd3se05UZtRWl/de9i6yJPwVpFh0lMsyxIfP3x0mn/Tpyn+/PKn7dfcEnF/a9Sjl1JIqNJqKrtI36nH1Za24fme64P+v/+//nf4nr+WvrkCHwi4gFNIDeqpzVOapPgj+QM/fvxo8GSu4YY0JqcGuOQwRTOUfA3XcQnQAlfXY6v/7aos3/B++L7vNh1C2B0YSef4nm819LhwgsH9Inl5tCOFG3IZ7fFxjO1tPa7nZKIMzOV24TUVma2OIKcqUKzfCABMVx/mMLCOnjYaMLzhBAJ24W87dxvca60xmUygtcHT0xOUUsjSzGnaAetNEGE4GqIsbZvHsihd/+/6sQUXl7lPPS4Coy0vVXDRsLXGGOSF1f0MgsBu0qv+4YRjeHvtaPM27LPptHmRQuL29taNuziOsVwuYYzB3d0dkiRxyiNdAYOdi0IIxFEMP/ABVFH6okbN2LFW7HPEydeJ4xh3d3f4+vUrACvNx5jtZhLHMVZV0UmX/YjzncLqRnJjd8VP0yfLL0jTzqQZTwFV4b5HR4KiGFRN1fidXgsAUzXym8nUGGtEozBCGIZIkgTJyupi+oGPOIrXb90y0a9xXHYdXdISfAkQn3XjGo2BMdot7o5nWK0dDNiIGtqPNQvX6sem4j1agPMsx8PDw5qPVH1Pnueu+Iuxqlc5twtf6ZeuCICI7lrrnl/bIQguwARbd7LhrcgSW3PgSN7tzQoeTeWccobReIS8yPHw+OA2Kr/+8itKZat6id7TJZAkDcnQZFnmUr/nQGnrLGdZhh8PP/D7H7+DwX6XgU2pl0V5FbbxMoUmtR016Wtds0PYANte7fqzQwrpJn+e250qYwzc406KiBaaUwb6JTTUDAyEEAijEEEQYDabYbFcQCubeguCoI+IvAIalbA1Oh3wc22q6Ppow6hMXcjd8gnJGG5EA1h7nFd91ncUoHC+jiwqpeF5PoajIZarJXRSFU9pOwcoVUyOqFJW9FhKCc444ii2kkFVEVaRFzY9id4x7ALIQRdCOGHzenRaClsQYWCFok+JhrsiJOoodIwMQA1C2vMLwxBhEKIoCvz48cOlifMiR1BWfO6y7ERBDMGtF2EI3/exXC6RZZmVW7vA+m7lZxL8+cefUErh/u4etzc2mpqkCfIidwGXLuMihSa0wxFMAHyz72GXF4ZtOwRa5Izunh7fa4B2pUEYIAiCxiCmVj6r5QqL5QLL5fIo3sglHWzaiYVB6BbDuhwHLXgk09FjPy7SxeeSFcJdqjbegnpkz2ZMDAw0jGHgNe0zivgBgOEkJ2KxbYFoRwzzPIdSGqPhCGVR4svXL9BqbWOFEG58O2dCG9cmjTZHUkp40oMU0vZaVuXBWmw9Xg5aW41PL/YwGAwQhmFjXHDGnZ7lKllhOp26jfprw/d8cMFtByNj9QnzPHd23WgryURKEO3x/aaSNDU+odEGaZJu0DVOPS5g52JZlpjOplZmSivMF3OUpc2cEkeUM95pObSLRApp0N7e3SKKInz79g1JksCTniPMdhGUeiFoaGc8fd+3KfAaZ/K9wJMegiDAIB4gCIKN51fkBTzPdq1J03SvU0gLDkVX3EZBNx23UyaJgUEURRiNRpjOpk6wmuRopCcdjYFSZ+683lnkdxvawt4MNhL23LN47t5d9N7W15ADHMR9Ds5J0ZEt3MLG60ClIUfnyN3vnK5ci6tsP7+Fs1SLDlGUkDFmBW8rGsdwaKOFFPVrRxjrDiVndvHL0swS66UEFxzD4dD11i2KYmMz1eN1wflad1II4TiitEmTQjaKkJaLJQq2u2jOySFV72/YYDzDJ3xm0661RhAGGE/GNnX88GAd1lLZLiG+B874zm4gddvy2hk42pwtF0vkXg4D4wIfVIHs6FFHnJfLkGAdSQWAr1+/Om4hZ9xpl9LPhK5pgV7EKWS8iiz51pFYRItqd9vNlmj7QCRs2r3ZF7sd7bwkjDFWiLhypDzPa1b5CuHaBNH7t4HEPh0hv85NNIDm2k2kU+8tVWHmRe76bzu+P2eObN9XYm5HPeW4LUK4IRC+iy9o1n//7D3D6440LTJ2QWkS1J8fb+tqZKAZMWwv3i4CU6WF4yjeoOlsO0/3TVVRWJ7nYJwhTVKEkRVHLsvStShVpernyhuAgTm9vMXCrp2M2YiSgXEOfRzFe+k6ztEgylPN5tadfsYYOHZEq57TntcaYRDC8zw8Pj463VrGGKIoQhiEWK6WLkrdDii89WacCndKVbp2vIEf2Ip9o188gvfW138ILuMUMgbp2QbQnudBcLvbAeD4K4QuKZxvBbMOhVKqIXT5XgylMZYoX5QFsAJSnq5fh128KIJI2OYIkGyCL3wX9WjIb3C2NkAau43UHlC1O7UJ00o7R9H3fJRF5RRWGoXvrYL8EJDwN9CM5pJT71pA1aJebdV/+wu4Y9Sjdc9F515zXm10tKmd27PnwWoOIVjjeu1Y38S+YoC280iV/HS8Zis8W+WsjYYnbIpxubK0jbI8jMzvzkXbfy8XS0hPuh6wQggnmFwWZWezOz8las0f8jzfcAqNsdqrvufvlCMiGheDjTa2NwXuOyonUyu9FlY/AsYYJGmCp8cnzKYzqwNbddgZDocIw9BxDH3ff7M09z6QDWNgyNIMxhgnvH0qDllTnD/R8RqFi3AKGZhrzcMYg+d5mIwnkJ7EYrGw4e4dKcauRBWIR+dJ68zWHdn34hAC6/tgf6hFMGqLYD0N/BwojUWk/Pp9dRGRE8YALZzz+dyR7YmQTen/oixcH8v3BOKu0LMikNPhnm/1WhAEDYe5/tk6Zw6oOYVVVMn3fEhP2sWh4AfMlWOe9Zb37hl2DC+9eTNVZrgmQVNBKw3peS5KQ2d08jeZmuRTRV/RWqMoC0gpMRwMkSTJ0dmY+uauKAoUeQE/8F3aUnCBUpQurey4kB2x0z8lDKz0V3WLiY7FGAMzDOBwhSa7ovpufsLAY2uJorocEaG++TiWU8oYw3w+R5qkdmNf0U0CP0AURSjKAnmRd56nSsoZ8/kcbMk27tEpxyM0pGuq51DntG88v45NrYtECrWxi0MYWILsp0+fXNpwNBzhjz//wHQ6Xcs01PCWDlfbsaHzL8ri3RYm1Em3gR8gHsSNCl6KLnDOkSbps8fL87yRgi6KwnJkarslxhmMaqY3DoWTcaicmFKVVn+KwarIl82oR5d3aJcCOYVCrqMKnHMXEQrDcO/nt0W4XJrZWPV+I+2CEka2kq8oChuBeDb92Pzd84+jzePb/YHnFri9XKo9fCv7u3Wfd/vvdbWxVV1I8PnzZywWC8AYtAUZ14cl5/uwc6wX8hlj24f5VSXybD5DlmVbP7MPjgpSifOXha0UFULAkx7CMITney617FQG9Nrx6HFBED+V2areKIpscKJ6nSrJPd9zklv7bGVRFG6O06Z4IyNXi07uOk4b7r1gjWYGjDGMR2M7JmczLBYLW/xkuq3HB1SbXrXWNz31fBufI1pU7ZjKqM3obUdxEaeQKlXLsnRcLqVUo4JVSusIUFl218CYHegUWn/P6RNjDDzpIYoijMfjRmSJ0o1FWaz5Lc9UibarKeuvn4ptKX0G5rhSSinLHSnLqzBOlwQR1aWUTuaCJE5OlUMg5wTAOmoMkqLhYGzd6rLxudaLXZr5u3b3Rx2jGoeLxQL39/cIfP8kRw3AznFqjGmkuktVIggCjIYjrFars1J0dWfYyYhU2R76Qyll6ilO/LTeObwgqqh8GIQYj8a2uAjrzjfUO3dplgc5cvXIfuNZET3kxEheWyBeSgnBBYbDIXzfx2w2s+Ox2pS/RzhbaWpKLB2PnNZxslNIA1Jr7aIPRVFgPp9jsViAMYab2xsMh0MAlXo/4xvOQWcWawNnEN+zQwisQ+t5kTsFdvc7xmwkQXqWq3doRNVsRqBoPFxqDHBhNdniOMZivrB81spxPVd24JrgeZ6tvq6cQsDOvyRJoEqFyc2k8f5GQcO5Gza23wBuOImvuEE8ZBE9BcZY+ZflYonBMEaSJmCmOd6e4xRuO49m9HL9jMqyRBzHGI6GeHx6XBdZnQFyFLTWrhq5LEu36ItQQCrpNvy0cX5v1IyXgEvpM5vSXywX6/FibCYliiJEYeQi8XvHcm0sOC4w1lxYBrZ1A/fsee5IW4/GI9ze3mK5XGK5XFpnsOLAds3mvmQhXD1TQdSaIAxcyr2Tfs8WnO4UVhVTjDMMBgNEUYQ0TfHw+IA0Tdc8JQOnwl6o7vae1UbDqNpDuyLP/iVQqhLL5dLqKyntjIgnPdze3drFSdnIwXMTzcleYHck5JTUcf29nHNEYYQ4jgEDV/0Og5/OIXT9ULG+b5RiqhPRiRNGFdi0oFAVK/3bpZb47uIIR/1o1JaYmsOyTi3Vx8I2yZQ6jrMH+58hA3NtGQ9CIzN9/GJRvzbq5hRGAYaDIebzJUhi5KCFvPp9/X6seYUchuYZMy6q5/s2C7NarZ6N1h8K4rIpraBytXYMq+IF37etwah9XlmsbQBFu3bx3npsh3vmDFglKyRJ0thcSSkhheW7H9K/ncZH49ioNuJ8M6LfmK875li90MzZAmYpRh/uP8APfHz5+sVFrR0XtWNZGiGF2+i07RvJlpHc06FD2N2TGtdeCgkhBT7cf4DWGovFwqX9aaPeVRztFNb5W0IIRFGEm5sbSGEFjUnOpP7+UpVOfLOOLg2WjcXqHRs12v07AVLG3TPngrt2S6pUbjHdt6iSZlWdQ+gizZSO2uEwHgJKd8WDGNKz47Aoi0o/rltG6VxQhNVVqVaajJTqY4whz3IX0akbKnIWi7wAD9eOIxPV/WkFfUzTA9woOGkvFNsc+81Fofksjn82p3MKjzjUzg+0r5F+pgr4p6cp7u/voUpbpVkUxcb93/Z5V9m8hXdkHcL1Ys6YbacVRVZOQ3CxYVv3XsVzEVNWnWt1umQHALspFFJAepbjpjzlxhpVolKUqHcOD0M96wZds5NUEAIDLriTDjpkI0X9kmlccWZT0FLIRn/f3RzaLecJK3NDn/E8Dx8/fsRgMMB8NsdsOrMFaOb5TdBbwfd8jEajRnEdYMcpOW2r1QqL+eK4jCFrpo2JcjUcDpHlWYPbTRvyrgbIjnYK6wMWzDZ89n0fSZJguVy6HaPv+/CkZw1jfnjHix7dAe0IS5RutxoEATzpIc3So3tbknEix4ZeOyddTzuvMAwhuECapFbDrVQ/Z2qr2qFzziE9G8EhQ0+cMOLytPtWE8qyhKc9xzfcapyeSQPvP8H6cUy3iIRnor3Q1aN7SilMp1NorfH502dwwW11IznwlczMrmj5Vp5s+73Vr20KVyGKIiuY+4Imts5BozEmpY2E+IGtPi+KAjrVzmbUncOuLn5dgos0bZlzVBVelMVBzn87KEM4J/tF63q9peXd3R3u7u5QFAV+/+N3pFl6ctvT1wLjzMmhNTJNzMqYUU3BcrE8/JhsLQOktXZFQlTs4/s+OOO28xa6PyfOLjThnIMzjtlihuVy6Urnfc+2Q0vT1Hng9d1DF3cRPTahjXb6f0IIBH5gJUiWpaMFAIdHBMigcFF1Min0WdEEmpC+76NUtp0QjTlKHf9MMDDwPM9xVRhja225KjpDzmDdyagbIarI9qQHT3quGGfr99HrLU7oTrTTt1SItL6AnwouElNpClKHHyEEbm5ucHd3hzRNGyn8XY7hoTAwgF73OKYoxNYq0wuBorCuB68qUZSFUxOQUjoxbFWudSw549DYXARPoYu8V/i+lQxaJau9c/VQnBOlchFjz8NwOITSCt++f8N8Nu90VJic2iIvMJ1ON+Yg5xxRFGEynkBI8SztpY08z+F7PqIwwsePH1Gq0gYqpIDgAr/+9quLQs7n850dX7qAk51CY4z1qJdL/PHHH+uFuIpikJfsRCHNeTuVlwY5rM7AvtNik7qxdj03mXKcvSiKkOc5kiSx0j2tXem2SErjZ87gez4YZ05Y+hzQ5E2SBACchIZpOyNXhDrJnMjaggt4vueKSBgqZ1CVbqEgEdm6Xt+2tGRRFsjz3EoD7YgmutQf+YR1539rWrBFOHSFEe337Ust74e5oJNf/+46Cd+dXv3ftffvSrfV08FKKTw+PkIphdFo5Do9ZHmGJEmcTBN9tn2s+vdZmyQghLSadYCLKFFhXBiEVqrE7ObtHoN9hQhEG6D7UBal3TTqSjTe96GldoUoRVEAGih1xXGjwjS2fWy+V9THIgVaiLNHagrL5RJFXmw4dc/a3IoLygVfC8+f0M6tOkEAdn18eHjA0+MT5ou563N8ahHLi6OaM0pZeaU2fQOw1zQYDFwWtE2faRyudd+oQEtKibv7OwB2bhD96vbmFlprDAdDFHnx8ziF7ciD0gqr1Qqr5coNBFMaDAYDxHEMA9t304mg1jgxXQOdk+/50EYjy7JOnudroO5gcFgphOFoiJubG3DO8fj46PSygOOeJxFwVanOrpqk71VKIVkl6zHY4dD8IaCuBAYGTFfC8EHodAeJW1QvYNhm5PahyAvkYu2c0Gcbz7IWHTwsIrzpFO69zmfGzWYq1TqGl4Dj/wDOiabCOAANMWH3/h0O4bYMiFIKT09PWCwWiOMYNzc3zqGn9Gv9/fXjkdNNCyw5hfXvM7rik4q1bqgxBoYdyavcdT3PFBy48+b2NSpsoEgoFxye70F6ln9cKus8ZllmHZ9679feMWxAKw0IIAoj3N7cIggCKxidWsrOsfdKCLuhBNZFf6dW4dbFmKdP08bv3HrQQa+QggQk0s4Ys+oZtXtAc3Ir37J1Se1rJHtN/57P5nh6ekJRFnbeCyvPNxgMXJasqziZU7hhIKsfOecYDUcYDAaYzmaOZ1BvGddl+L4PrXWnPfnXQr1Tzd3tHTzPw2w+wypZNaRejjyo261d0nmrR7WuHcaG1eFLy9eiiF5ZlLaIRJUnO4OA5c+UygoTSynxXOVqW5vsubN3YAabYtPX/ZDq472eOq5nFog/SFWgRGkIgsBVHvq+v9Uh3PY8SQeSFiI6RpImGA6GmxGNNzaxWmlXvRmEAXzfh898W5hW6dhuozX0qFBx8kfDEeI4RpZltsL8xEg58d1ISgh4vwVAxD8nnqYDW88rGrvn+CrL5RJP0ycUeWG531zgw8cPAHZsvjv0PC4iXl1HHMcYT8ZgjGE2myFLs6tJxTJmW34dU8n3s8FFIqo01GAwwORmAs/zbIXZzFaYGX3a7l6VamfU5exzRyv606GJdsw1SykxGo7ccyhK2+OWromiQhThOkVKhRnmigY833OO3yGt4nYR2atXqi+hdPJzTmG3N4m7sC1C2KjMbkUbZrOZ4zF5nrcWtd1TuOJgGOr3iXEGKSTyPIf4VXTCESTUu21orWFS43i/nHFHPyFe63u2tbsQxzHu7+9d7+DpdGq7R7Hj7EgdWuu+KUO1gfN932ntEoQUYGDI8uzo1pEA1godFWiDp5TdCEkpXSEL2XJ3Xh0rxjvKKdwmmUBNuwUXYJy5KOF8Mcd0+uR4Z12MELZ5GRQ1oX+TnMT23Xv3rudSEHwdCpeeJZBPn6Z4eLAalHVZgmNRqtLpQV16XDDGXEsu3/Pdd9R//xYgfqaGdpyewA82+HyerPiCnDnKRf0PjU36j4597H10hT6skq6oKuUotVdH3encVSywFQbY5qlsnucxz+Rlnp/jC6KWNm07WgY2f137TOPManaCnHbqXVyvTgawfp4Ho+UUVt9VliWyPMNoNIL35CFD1uD71d9/DE6dJ3UlAeJn089a2yIYadZamsYYR4WAeb6/73uB79uWsWmaYr6YY7FcoCzLDcfjUNT7WF/6vpJWsVIKWZYh8IOLHv+SYMxmW2bTGVbLVYM6I6XEYDgAZ9xp6jY++wxXkjrQaKORJImlS9Qk0aSUVlYoLzrf6eV0nUICW/fQHEQDjEYjqFJhNps5UmxXwRm3sgq+rZT2pOf4XOPx2BmsoigcqZvQVUf3XBDXhyJGSZLg27dvmFVUAG00mG4uUMfgnMq3fahLJnB0i7NBjgZnHJppxwv0fd/yTTzpokdlWaLMW2MN66KZbdIVR0dF2fo503cC1aK8r3E7vX5Q6u/8udEeWy9lSpxDaGqR5hq/EDhuN193DoHNMX9Kgc3G+VbFe1RFTuT418Bm68LdRQv117TRKEq70RbcOoauJWWe2014ffF9p85hmqb48fDD0kWK3FERtDnNqTt+E3IYSN6FxjeNw66u+QzMFebVN3FA1XM6jhy9aeMa2Oa4b/y6uu48z/H0+GS7R6kqK6aNazGa5ZkLinQVF0kfU0rk5uYGcRxjldiy664LB0dx1Agl1x+W9CyBO0kSJxja5Wu5JOg6tbbV5fP53A3wdoi8KzAw4OA2AleF7Y/VUXwpaKMhmHDzhKIovufD8z1wxpEkyZp3y5mrPH4JtJ+bUlaIXAqJTG0WWG1zAnc5hscWjxx13tjfmUa31beP+G7nGNayAs1FwPZ4BrARAaRFsf4aLeTt76j/XT+v/ef2vEPMeBWNfmNtzl1jp/6zu1/KRm7CKHSp0iKvRbU6llZ7LZCEkRvvpnt0GMA+yzRNncOzLUrduXWTCslac46aMpDwP4Cj5J2IJ6uUwo+HHyjywkpEce4aDEhpGyu4bi/V/WJYt3ztwjM+2ymkarPxeIzJZIKiLFxTbHIiurZzoBQcGSA61zCwuwWtNbI0AxjcAOnUwH5NVITbekq5S8+zISlgNAIZQEgrYg2czsF5CTBunULO150FiqKwfWbVdv2x1xh3lMaL4qjb4/yZgphLLpwb7frQjCLuGlP13x16L58bo5tBi3VU3P7euAWFIsldh1sADbBarVxXHh7YIqh6xXIXFsrXAjkINCZIb7WT96A6pbu7O0RhhKfpk7O767ecVw3/WiCtTWp8cMjtblNriD6xWq2Q5znCIHQyQOQU7pVhe8a+vRbOdgrJwRJCIM9zy4GgPn+6A1e4Ba6QQjOkqR3Enu/ZSr7q4c5mMwDrdk31FlU/M3bxxhoRlDMcB8aY2ymdc0+3LaLGGDDOGvIA9J0v7RiSrhh9LekLUmso6k1MVIXVctW4Ds54IzKyrZn8rkgZfQ+hHi069LrL0vaxpc+0ebTr49AOe/3z+g8A8Ip6Z50To1vXcERv4k0OMwC2JxLWOK9NsD07/3akb/ubqs8bjaYFN7Xrss+QMwblFBcokmjWH2+f297zRqOIm8Zavcq5/gja0cKXpFPsG3v0+/0HgHN+SN82YAHyLLfKFVDrvunPRIrbeOuo6akwxgAa7rmecu11aKNddPvcTZ8rRKzWUCEEwiDEb7/95hweUjagwo4ugmgzQgpEYYTBYICiKKze8oHpXRr7dWUVuj+uh3jVdci2vlTO32jY6C0R1rfERdLHxhgsF0tkaWbbn1W9MLelULqEOj9LSrke8Nps7dPc5Wu5FPbt7Oj1c3etRPA9p/LQOVwtI0dt3+qhf1fo8UKLhDHGifOSYaDzIM6gFFafLssyzOdzVwjTuKYan0qw85umHzNetbZ8Lyoc2+X8mw3Hq/mz+8xO5++5auTaO1tz7tk06ovutOsH3/ZF9Nr67/X9Y2CMHEkAfNtJ7l+seXuDwFhnF9xjQfdJKdtH2fM8+IEVuE/TFAa2UcIVBJzOhrOt1V9tp/tYUJcb6UvnfJ+zsafPcmGdnqKwQvhKKddqk8Shu7xeMsYgpO3QNZlMHFUsy7Kjzntb0ARYy9sEQYDb21sYbTBbzJDl3Ze6O9spNKYSsU5W1muuKm5eqqDg0iCeVxRGG69fw/m/Oi6w8AaBrVBbrVYnfP16sa334aTfSSmtE+ZJ16LvVIL2wefErBAqY8w5gNKTtvl5RahfrpaOP7LNIbw0jh272miURWm19Jho7JYPmcuN58AY4JzD/RyzY/HcYraXc7hnT7C1irv2zzrH0NmG6ve02XBR1SoyqMvtX7jb2T4M7THfJbR5WMdsxJxzWCrH6ab7UqDobObp4qC9xQVAqegwDGG0wSo53ubWQfq9vm81VMMgdAUnURRhuVwCqhLg5sfx8l4TxOmOoxiTyQRgVvczz/KjxtmudUVwAS44RqMRPn36hNlshoeHB9sUgzOY8jgu9mviIpFCEnumNDLQUQ5EC7Sj8T0ffrBeqOncrzX90HX4ng+w05zCeqjd415DawpYy7pIIWGkgeKqUWH7UiDOSBAG1lAyKxmSZqmbG4wzl1Z4sR61JzpdVN2ojXairruO1S44qe+Wu2TczkJr87OPr7jrd6TKAADPZXD3cwq7b0tPRd0Rl9I6gmliVQ48z2tInJRF+a519s5BEATQ2sqlnLM2h1EI3/MRRiGiMLI87iBAGEaYTCYwxiDLMtfrO1klF7yKM8HQqASOoshq8PoeptMpsixzjTYuEaGNPNuRRivbEnC5XHY6pU64mHi1q1g9llPyxojCCEIKDAYD/PHHH7i7s30Lr8GpfQ3UuSPkWDWU4PeAxgLntrJLcIFSlYjiakd5JhhjiOLIGqdqsfB8DzDWCAZBgLIssVqtUOI8p5AcuTqfhq6NWidR54A0S2H0mnhc18N6aWyNeO1B3amjRZcI0o0IoSG6RZNjuM0ptN9dVeru4wC+Mtop2OeqlevYVpn8XDUz+DqSRzJOW7mwz9iardxSvpZ1oeO2I7ptm9y1qA3ND86takDgWy4hpSZpTjuSfpZbztc7EbzWRq/5aUc4KL7vY7WyVa5RFKEoCydcTWLKu1Cnjmz7TsYY7u/v8csvvzi7VpYljLbO4d/+9jcYbfD7H7/j3/7t3zbG7luNQaJblLpEEAa4v7/HIB7AD3wsl0ssFouNsdXmpW+7H07aq9Wxjdae33//HUEYYLFYVFxj3vmNzcU7mlwTpLAt3EajERaLRZNUbzYNeNcd3JcAFxxBECAKI8sdXS6t2OwxMHaHBr5OtVKjcOD0iGxRFJjP5shSG5IPwxBS2rRxqUpX1XuJiK9SCqUpnXHhjLvIhuevNQaJYH1toJSJ0QZ5kcOH3+jR6YpgzHrhaP/5qSKFLZxCJ2lUItNCvLXI5Liqaed8V2m7ujO+jWfbNWewDnJ6fN/fcFbaY8rzPReJ+pkdQ+L9RXHk2txl6eFctCS10UAhbcFdfVNKeqjP2URXjLnFGVosF/jHP/9hnRzBcX9/j5E/QrJK8OXPL2CcYblYQmvtModdQb04y/d9PD482qrpNN1oVQmcvuZTQUmapVgsF24jd+n2ri+Bi+kUXiOIeyY9ieX3ZuSKcdsK7L2DwUYkhsMhpCeR5dnBTiFFMojnRzwL6dmuBvEgXqvtq+cNVRtKKVsxlqXwfd9V+FKhEE30nRIAx8LACU3HUQzpWYmBJEk6v/vbB4pqEVSpkKPpGJLj0nZe6h0srtUOHAvGmt1PnuMYNrDLP3tm+HR9ITkHVLjwHJeLc+5oPj+zY0hzLo5j3Exu8Pj4eJRTaIxBHMeOuy24gJACAgJDNkReWKFwVaqjnUOjDRbzBeazOYwxGE/GuL29BWCd0e8/vlunS5tOOYTkDDJmpegeHx+xWq4shYnBdd85V11jFyjyvS2S3zVcPFLYrsLpMqSUiKMYDz8ebB9R2Z1B3BVorZHnOQyM5ekdQ8I1BvEgthW4Uro0qxQSqlRWTzBNHQeFWtQdCiGEi+jWq8epCi7P83W13JnVx0IISF/CD2wLKmC9MHVtrJ+r12eMcY6hh3W3DMYZoJlLawHNlPFLGdQePy8441bQHcxV8LdRH1cUVQSwEd25VpDqAM2pwA9cFkIIcbR9CcMQN5Mbq7mrmkLriIAsz2z0McucTmp9Tm+Do8yYtXi77/u4vbl1RSzGGIRh6GRdpJQvzuU+BtRqUWnlHMJ6luMSoKi88ITjLiqlUBblVTiEwJlO4bYLm0wmuL29xffv3/Hw8GB7/nWUWJmsEvxj9Q8AFT8tsuK9qtzUWHxOJ6rOM7t21K9TCOEEOA2Mjawq6Vq1kdHZhdVqhSCwXUbSNMXHjx+RI0de5Fg8LhD4geOyHXv/GFhDST/wA3jSc2X/9fM61iGkNHGe57Yv5mCAIAhcj0+SYOginiNJt7l0GzQJvhbOJc6X+yM4RFXRSFWNUkon5bCRumzN/TddxNvn1grbHcMxtMezf+3jGLY3yTvnyjMmstHWsLr3XPNGUdC1cQo55/BD2+qR2o8RL7eN+tgiEfhSlZ1vpXooOLM9hLXW1qFi0gndCyEgPSspQ9JW+6KkSik8Pj1isVxACGEpLp6HoihcVkMr7VKZzzmEdTDGIIWEkAJKKfiB74r98jx3BSaMs05Wi7sofuXgAs052VBQOAIbVfdKYzKe4F/+5V/w7//x75jP542N8zH3/LVx0UITBobADzAcDK3mT5rt7NTQRYxGI+sIMEt23iUp8TODMWaLNQAMh0OMx2MopZxT9PHjR9sLuijx8PCAtEz3TiDSsBJCbDUS1Ff6EJ7L9hO23FCqrqN2Q3Qtp449ImV7nocwDCG4cJHHOhH7Wsb2MXCOjLYbHYoMcMbBBWv4VlmWuefXw+LSLck2Ck3qHML6H87A9PVwChlb68Nqra3ju0eOpc4xpLZkSinX9eNaYWBl3cIwxGg4QhDaTXQURpaz9+Eek3ICVSo8TZ+QF/nOYymtYJRxc1IIgUE8cPe4LKyOIKWOj42S6aqgBADu7+7h+z7m8zmCIIDv+85ZPYUO9DOBIqmlWvPQnVSV6q5DCFyiowmaWnFc2J2NEJbHcA3ESsAanIeHBxhjJ1RZlp01pi8NMiaT8QS3d7dIVgmEFNBaYzAYwPd8a1i0Qvn9eYegLEvbrSAKGwbImKoQ5ESHkLgunvRslV1RoCiLs+UEgHWkMAxsJIwiGZzZiBkYwMx63F9rpLi9M25EtBgcP4gxZiNpylabOFkgz0OWZS6i+B6xj2PYrkrchXNspHMIr4zXSU4hDFDq0t7DPZWxQNMxpPTktbfCo42m1hpBGODm5sbpCyqlnMQVPVvqEb0NlIqubxZ833eb3DzPN6JUxxZVKGUd2E+fPkEphdVqhSiO3HHeu0MIWD8oiiPA2GrwOI5dISKMXTtcYevP1tGEGrGTYQLgdm+kCbRtAHYB7YE7n83BOXf6WO2CivrDO6ftUJdBOxni7cymM3z7/s1NdCFs0cnNzc1BToCUElprSCExHA7X4fNqt3RyhLCC4MKlWcqibFbbnTHUKO3ie3a3R2kRKeWLtg3rFNja4XFpF61RdwrbnMpzorPXhLe+zvqCck1wUeeKjlDnEh7KS6X3SCnhSc+lQ685Wm2MQZEXrtXaYrFAnueOC+37Pj5/+mxF8fcEK0gHVUjh1jGnImBwFGd7G6S0LsPtzS244JjP5s5JTNPU8ROvBTTmLs4trHFfqY0eVZGvVitXndxFnOwU0i4kjmIMh0NwYZ2pwWCAKIowGo3ge3aH8vD4gDRNXQpxnzF9rQG1TW5GetKlBCnsWz+vhnPbMe/+paCUwnK5dJVTxHEZDAaHXb9Z92oVXGCxXGA4HNr7eQEDEkURoijC9GmKNE0RD2J73lptPLNDJzxjlrNEWlNGG8ubYbs7SFwiOvlaqC8qJNTajhY4A8ks9841fmeAqfVlJn1GWuzrx9j63W/JMXzm+ded/eecra0LCHEM9bqP8jkdPp77bpLOqp00gO6mi4GmQxdFNrpEtJJjzpv4dUEYwMA4buE12mTG1r3RqSvYarWyQtPappZvbm5QqnLdB3rfpoTZaKIQAuPxGGmaIgxD2zpwy1w/Bpxz3N7e4vPnz3iaPmE2n8GTnuM5Ms6AKyoKJ6e7rkN6Cfjemms5HA0RxzGKvECpSvzxxx8/n1PoQtNgGAwG+Msvf7EFCVWUTQiBT/6nRgXo129fO5WS3UVmNjBWiobVQvG1xf5aKojOwT6H1/GAwDYqqrZ/wN6/8WjsKtHqu7NzwFB1DalER4UUbid70LntgOBi3ZmnfQx65Obto0WvgnZnD8bAaiLeFPX5WefCLux79vWI10Yv2y0bh339xrd/wfp71i9dlsf4UiC9Uk96Vsy+XBeZHZv+NjBOL1Srl+9a9JpwY6viTJM9UqV6lqpCXOgoimBgkKWZU44QXJwVLaTiwuVyiaenJxRFgSiyLWKjMMJ8Pj/52K8NosZ4vgem2UUljsbjMbS290lphcV8Ac+3gQZao7qKo8+OnEEyYvP5HOV/lo4Y++HjBwR+gB8PPzCbzWC0FRvlzAr+Hm0AXwDkmDYI2vWigWohdFGM1sL402OLcDfBhcWr3Wg9QrT1UNpgMBrA8zwrqmrWz//sqAmzfEUqZiK5G621lVo4cqFxkVApDpaCaHPxrg20U95bJcvXHBhajK6Nv3YJtPmwO6+/Zi9orFM0bNdnjhk/9XnTjs52ZdO9C7SJIGFlsrFEQToKZt0tqe4QXlP68jnUo4jGGOuUVVkbGjPtZ05KDHEcI01TrFYreJ4V/rayUqefD+cci+UCWW55xHEcYzQauarpawHDOlodRRFms9nFnELGGCY3EyhtC4NUaQstb+9uEQSB46R31ac4yWWtO3ZpmiJJEnDB4X/ybUqw6nm4WCxcCJw+B6BRXfYWDiKdvxACnm/755KxcjwqY5BnOZRWyLPNaq+feUEkY029ibXWDUeRDBRV+u67F0IIR7LNssylD1317okzgyoVidNGvJlSWeI5RShpI+I+s+eaAWtgSRbDaOM6eLQ/z8Bsl4/6z1fmGB5976vimvbnyJk+BXs3FEfez2cjt/Wvale5VoUh7q2t33fx0bbvnWlfQwfoDI0sS1VIIoVcc4DPuLEbc5ZbObFrhTE2gAKGhoPCObepSAPXsq7xudZ8ZIzBD3xwzjGbzaydpv/OHMhaa5sGrWg14/EYUkos5gvbxeRSjQJeAPUiHBgbgb29uUUUR1itVsjz3G1229SMQ+aSNlYHkTqAPT49IlklUFq5Ht4UHe8yjnIK25WWTkqAs6opdujaFQkptkaE2ob7LZwrMp5+4GM8GiOMrPgmqeW792mD5WqJL1++uNd+ZmfQwdg0wR9//rHBlZPC9iElw/AcgiBw0eJ6azuq4i1V8xgHR/Vqjho5JCRvU6+4q3NYnzs2pbGEEOCMIysyZ0DA0HQi2rSCDkTAn0N7QXDFClv4tdvS5uTE1x1gMp4UrXnr4ov9z7hh5Zue3taf28c//xwvgTqtxVExaie7a7y/te1iYOByrXlZ6FYh35FE/zqFgVKs9S4db329x6JUJR6fHt0mi+R6OOMIw9AGKCo6Vn1stuccZ1ZXdjFfoCgKCCkQ+AGyPNtqs4+5T268Kfud89nciWAvl8vO3vO6SgrpsAK2Stj3fMsfLyp6E2euy9ahoPnneR4+f/6MPM8xm81QlLbamGoUlFZIkmQrF7grODm53U4jUdk1mOU9qFJ1WqPQVcHWdj5155Uz7vT6KF1+DZydS8Glu6oFiFISo9EIggvMV/NnU8cAXDcUrbSVjomjtTN4IftBKWljDAwz62e1h8d1+MEvc44/Cxp8uQtW610DGuOIbfKLD45StnHsGKs5hPWf69SMrkJKafXbirVzcuoYavBaSbewVD+Nviw5h0FoU45U3Qs8E+VnQJqkrtBuMBjY8VqpgVyyuGu1WmG5WrosW1fX+zoPVwrpigkZs7x03/dhYuOctrIoHa3sEFBRGRXZzudzZGnmslYUTMnzvKFTuK116FvjdKew9vAFF074OctsdKVUpSPFdnXhWC6XLrKUZ7kT5QQqj/8vn9+lU6CNXk8GZtMXZVnCD3wMR0MwzpBmqTNa+wxBnud2c6CNrVLnHEVZuFD9peCiJRobC/BB37PtEgwaKeL3hF2FWPS7Ls/rl4C91no+ufXjOfeD4Tiel6lxCWnhupJHQfq1aZpehP+ojYZgwhXAFaIAyjOfR4fAYLn6jDPr6FXZjH3ZNmMM8jx3qdIojNbtSi/stBEfmcFG17qqVUrZwTAKMRlPrEA4GKI4guACd+IOWmnkRY5vX79hUSyO2mDRpowkheaL+boLGLcOoZTSFZ6sT+wFLvZMXKQMJo5jVzJfpLYayWjT4OcRurSTpV2CUjayWU8B1vs8/kzE5UNR373QroqEnJMkcSKojQpLbD5fY4zTEcvyDNlD5pzMdhXWOUacDGU9WlJ3bM848EFocwwvddyXRGOs02s1usC+HWxjXrN1xuCSi84p4+HVIhUVv7L+81GRwy3HO/ytzeISoOkEdcnG1sEYc235VKnAZKtYqX27DrwMss9UkFEWJfIi76yD8hxcMSdjCKMQQRggSzMsV8uD1qK6HeSMY7FYQCmFJE2gSrXWLcQFUuzG3n/q79umYHUNgguMxiOEQYjVamULFY3lXHLBEXsxwih0fPpDQVnHNE3x9evXddCkkmOL4ghSNGlXXYwSAhdwCqkptu/7eHx8RFmWdmfDmBMWrZNmu7R7Y7DnGASBrWSrTRbP89aGvnpu27hX7wFCCEShDYsrpTCfz5Fn65ZvDbS4diSlwKUllteN2iWjhdscwFd9Puy4xfgt0iy7Kozb533IfSMnpF2F/PPOif2RwotGDp+B27yy5jOlSvJ2BK5Tz4RhLVxv9FFC8Ls4ko4fVmmocs47sek6FXRdnvRwd3sHzjh+PP7AarUCFdgdegxtdEMmxvO8iwY5aPPDuU2ddrmnL2cceWHbriZJgj///NN1XJNCYjAcYDKZ2OLEE+Yv3YvZbOYik1TQSpJsaZaiKAo7R7t5m853CqPIqnUvl0s8PDwgiqLmIoHuivpqozGejDEej5FlVsuJ0C6q6eglvApI7kUIgfls7iqqupqiuTj/80iHr0ePVwWr/d3RhWYr2o71mSDNQi741UYJCQbGdi/hHPP5HKtkZdUWzHFtY196c0LZIlo7t6kTdAFUYELQxmauSL3CeKbhSDN+mPPd/g4CF9xxFYfDIXzfx3Q2dY79OVHC59aic+//RdLHSZJgsbSVToPBAACuInrgebbMn3iF7XOupyG7ONBfBcbu7CnUnuWZ0ye8JE66x6Y5AerFT6eQ93e93tXx2+N6cO4Y2ucIXNuGZZs02SVAsmJS2krka7XZxhgnXfLw+IAkqdK+nF+Up3+JdY1z7igBbc5x18E5t+oUbB3Vo44ywCYd5BgIIVDkhW0LOxgCAGazma254MwVDJ2C587l3Ht/lFPYHozGGKxWK9fkeTgaYjKZQGuNUpWdrj4GrDP4+PSI2XzmiMrG2JZmcRxjOBpaEeRK9PO9OgelKlEsC7Alcy3NDkGjOpJSlWaTD1WWpdMvy/N88/Nb0JbhACyVwfd9FEWx0bf62XPFmhNH4X0hxUEV1ifhDYZSO238lils+v7nnvGxEiUHSxptsWV7z80wYN+5bkgSGdR3Js/f6v1vYBt8VVOdjoEB9aNu9qXeRRd4S2itG1qljTHYinQe67SQTJoQVny+LXd1LSDblmWZ1S0062s7BFppSG/d2Un4ovF7Yey94ZwfXRzigiemspmc4fPnz1Clwrfv3wDYdpEaulOZpDrVKcsyOz6K0q1liinXmcmJg9fHXpsldYBjxjjDzc0NBoMBFsuFrR4nmscJCuLbCsq2OeDu3FpBk0NxdKSw/aDzPLeNuznHYDCwosfLFbI0W4sbd3Qnq5Rq8B2FsNqKcRy7IpQ0SxvyJu8NxBGhDh/HGFpjjJWwkWInz6lUJRaLhRWy5Wbj87sm37bJIKVEFNoip2OdQgCOS0JcxzAMG7pnF8VbTImOjeHnIgrHRhyO2UFvFMA98/NzqdmNAqvNb997bsc9HJoXNcfQ1BzDjhacGGOcE0JV0/XFkdqL1t+/cQ17LqmtRXdNPXjroHFMfGyt1s0DDpkTQRhgOBzC82xPYjoOHZvW6KKsNs9HZNrJiaJ7LbnE3d0d8izHjx8/LK0IptE0oAugjjlaazw8PLjghtswVdw/pW3RKd1vh41h+PzciuPYchQ5x2K+sMVVOCOK2qIx7Vwba/z6Q8dMHRdJH5P20XxuteuKsnBe8VWhKjbxAx+e77koaJcd25cG59y2MhqOkOUZptNpo4fxc4jjGJ7v7XQKjTEoixKLwtIPDjlmm2Tf/vvUR0U7YGqTRy2J6gLYPXqcgnMioj/T2NNKQ4RirZf3Ainkawc5KMPhEIwxLOYLa3MPHAZRFGE0HLmmDI1jVyn2mTfDw+NDw2E8BEpZx0Z6Ep7nwfd86+xrZXV9i3VP4S6BbHtRFMjSbEOD0Pftmk/BrHP5uVJKTCYTMMYwnU5t5fiWtPRJ10J8R7ZeCxv83LZDe+y5n3V2FajiK89tZQ8VIQDd263ugzG2LJ3SkLPpbP0gO7TreW2EQYi7uzvM5/NGJRtNtH33Jk1TFGWx3SlkwCAeOA0nA/Nsl5S6aK9LZbDav7F9zDW0F+vn0D5+zTEsy9IKnJq3S7f2+Plx6YhpF0Hnr5SynD8ukOc5hDzOKXnuO8gOdM0pOQoMLvPGOUeySo5qjVYUBVbJClluO414nud+R5Ww0rNUKSHFUT1/BReQnkQYhgjD0MkACSEQRZXsSlk1g6ikyBqX9kZOu1IKRVk4p5ibNYUBsPUFnvQwn89d95FzEIURbiY3yNIMD48PKPKiIVh9Khq1D+6v5s+vyilsw1Xr1B48VfNcS8Vm/QZyyeF5HgbxAIILZFl23cblAuB87SS7CVXvJ/yMY7hcLhvvFUJAKw0uOMIgRBzH6+ruLVnaDRmK2pgyxrYmjOPYLQhknIhbWJaljfbqLRXkex4tib36vu0hemgUs8vYxTFrpCRqTre7P2x3NGvDQb8gLs1JOiZat/ndDMeEtTjYxbaR++79rj/t97023ALYWghJy40qQevXtkHTOTJa44Ssr2Dd2QdSe4ijGKWyFax5kTsHTym1k9fNGEOe5y7DRRx5uiW+52M4GDZTp0eMDy44hsMhPn365BypKIzgez6iMMIqWYFzjr///e8oimLT4Ww939d6VsTJrNtAxphbh25ub6CNHZtlUR7F4dyGNE2xWC6wWq6wWCxcdfY5VCRj1h27qMahrhVL7wHWG8lTNpQXiRTWVc3phK4BbmBUApNCCEzGE3ieh+lsiizP3EO89p36qeDcptONsVE8T3rwPA9GW35hWZY7e0QaY6yILOONEn9VKgjUIgSmSQQmPCdnZGBcs3illHMCCVQ4RAZyA88MU9LYbDhK14xaeqH58h7eZrVQ7zMu9XtzDK/v2dO9cISsfW5HcQqBozYVxy54x0YKNygTza/GMQ7sS4KcwbqTmGUZfN+3G8SKs0zFDg0h9RbHsHpDEy0OInD9kVUhBOI4hhACWZ5BSIE4ipGLHFmeOTrTto042WlncwEordYBnNp6Rn+OcswMXCEmOfhpmrpfB36AIAjcM9g3h7Y+3xcE8eKBaqxwS2+6vb1FHMeYTqdWfxfr9omnoigLPDw8uPXRcHM2N518rHpRZP1328b8KRXmF3EKrxXG2NJ/z/Ns0/AgwHhsRSa/f/++bpB95UbmHHBuo6dhGOLjx4+4ubkBmO2t+f3H90Y6uQ2aVFEUIQgC15xdlcoaujg+69zImJWqRJZlG22cwiA8+bkx2BRUmqQIwsCSkI9Is/TYjks6jT2uB3UnoSgKSxnx5DrNWKtK7rFGFEYIQ9tJqixLPD4+4unpyVUl7wJp4+VF3ugc1e4ita2gYp+T6LpYaYPFYmGLS2p28bfffnOp6a5DcOH4l2VRYjab2TWKi7NEuOn+kLPMBb94saJz6Fubw3aE/hS8mFN4LY4U5xzSkwiCALe3t06mpl4ocw3XcWnQ8+Ocw/ds6lhKCcZtq6o4WldoL5fLncfxfR+TyQTxIEaWZs64ccExiAdI0mQjBH7MOcLYyCPxWTeiQTixSITZz+aF5T35frfbN3UFz6WRL61v2eP6QMVlgot1ha3eImFyTsHYFUNKy9kDrA3yfd923vIDCG77Ru/rYxxFEe7v7xFFNp1b5xQCaNJBWCti/kz0jmg4xhgkSYI0TRtOIXWrMdp0mnpFqWPARvWmT1Mkq8RJkHFYR+5U/p8xZvuYPuN829Sp9rEvNe7Pcgrr4XqlFDzPDlwq66bm3ZdofP4SoEnx4cMHRFGEPM/xNH1at6l5pzDGuJJ93/chPYnHR6vnqJV97cOHDxs7+/bABYA4smmG1WoFo02j6lApBSnkulqtNaa3NX5vT4z666q0TqGQAoKLjZTJsSCnk/o0UxuxS+AlF67nxm5d2f8Ym1ff6LW5hJfiFO7j9RkAZt+C9cy1NH5vANTHr2mNP2OA+vWYLVSG+o8bw+K4e9GYS6b5ecvR3pIaYgIAB2PC/eGMgbWLuvgLjrUdCz89N2pj5yhG1etFWUAbjTAIHedNKeVSn1xwnCXfcWUgmyulROAHCIMQaZZiNrMaupTFUqVq3PNtcy7LMqRZurZZynboUEphOBiiKC3XjzO+tsd0HgfY3DzP1/ZbSsdx9DwPUkpopaG0ejmN1xNQ59jRzwCwWq6QrBLbfq4s3LWe6xASLY06l+zzgYx5vrtJm3tLjnde5rYYktZArIt821SBje/cMbcuEilkYK4g4fbuFqpUeHp6cp1CugrBreNT5HYwLFdLzGazhoDyewQ5Q2EYYjweQwqJ74vveHp8Aucck5sJtLEC5c9FfmbzGdhiPQZ837cGRHpW9sUPbAppS8/WDdTL7isordwCs01Pct/gf+67aCJqpaFKawB/uoXqSDL/s4e7YMHJi2Yb2tfNWNNr3PgZ++/TJe8jY03vd+PYtcVtw/l8ZXt75HXX08hKqbXzwjmkkJDhOqVsjHH6cu8FUkjEgxhSSixXSywWC1CBH3XbUEo9WyS3XC5tJC9ZpzBhgPJDiTiObUHoCQOWcebsoFb2XIy249GTHqQnXRSzy4odDAxlYYsQHWfcAIaZ09eMGo7itx44hxoC+aYVjTxh3u96Pic7hY0cNoOrQhqPx0iTFNPptPMcES6sjM50OgVjDEVZ7A3Ldw00ELY93FMXVDJASilEUYTbm1sURYHZbIY0TREEgeOllGXpUgfbooRANT5qp0FFKcRTTJO00flmF6F+F2gBeY7vd+zCUi+wIO1NIcTV0CK6irZNaG8qrv3eUvahHdJ86eui+dfVhXhblJ2KIih44Hu+q/Ynu3HMvHX3/spQL2QjrnWpSiSJlaKh4gLpSaRZaqNwZncUjjHm+Gwk4u/7PqSwUkBlYe95WZQbDtBz91sIgcfHR6sqUfFDlbZZQs/3EAQBnp6e3DrSVbqIga0nkFLaAEdZVRzvS0WcAEpF07+B020BOdpOIo3mOrGvKi7judmsi3EKhRDwAx8M1rnSWsPzPZcS2LWYvmVqmYzPcrXc0HO6ZtQdtFMqqYSw6dc4jsE4w/Rxivl87viXUkjH5ds36bXRG8LPxlgtSKr2PrcVoioVStQ0vNop6C3ci0NhzLrhO6VEpJS9Y7gHuyKF7bTzT3v/3sIpMbhotPe1QPwzmmNFUSBJEwRBYKuT5eEtNR2q+/AiXYheEGSzScNxuVgiyzKrrFBVD0shDxbSz7IMwHqNY4zB8z34vo8stwLN27pT7bKV7jVjo4XU9UmVVpeYnE5Pera/b8edQsBmwm5vb7FKVnh8fASwO3p2MZyZUSC93fp5Ghin7qH0+cWQRzmFDR5RtbsR0lbweL7Na3ueh9FwZDlkxqDIC6zUCoyzrenkt5y8NLCNMZtVWR0GTVwq/qBUDABbPVaFwum99b+B/btBxphzCu/v7qGVxo+HH656mIpEACAvbJp9p2O/ZafPGIPv+45Inaapix6eQkxuOMBVYQyNS+K2nhRap/tWRQwNLIdDCgnDDYry+DZ6247/XtB2Bh3nrBY53MZ7ufT3Xgpb5xDb/vtDvrt5PNY8WGseka4npVYpgpAXeYNL2wXsuv/1cSCYLTYxsOmwJElQ5AWCcC1vQp/RWu9PnRp9VdkeYL1xD3zbnk56VgCaHDshBIQUtlNYlm4tqGscr84/M7ZQRSsN37PFclSo0n7v3nOs3U9y5jnjtjFB5fxNbiZ4mtrKaOK8dQn16+ScIwgC3N3dIUoiLBdLLJfLhpj6ruzXMd8nPYnffv0N88X8Yo5nURROL1gGlnrBOXfP5dz5f7YnNBwO8dtvvyEI7ASWnkSWZhgMbR/kx8dH/PnnnzujhW9pwC5VGfRWoHQJhcEJ2ui1mrw+7jqpMtAIg6fpk4sIUuulIAjgeR7SLH1e3HvLVwopEIaWXE6cDmB7eulY0OQQ3E7soijsbviMR+ycQ21c2qbH5fFSi/jbkd3pOy/j2B50f7q1Bj8LxpudR+ppVKWUpZaUJXzPRg1pfu/jfNHvrs22O45lmgIGzrEC4CqPy6K0OnpHzpWiKDAejzGejME5t/e1OLxVafs8nRC50S679vHDRwR+gNl8hrJYc0K7CpJaK8sSi8XCFc1cujCWMVvlTJvfc8dkfXyDr4M4WumLdGIBTnQKafJSiNgYg1Wyct0rkiRxQtDUmDtJkk5VI/0UYNvTdfXnU4/qHgJjjBVMFQJfv3617QuL3BHB4yhGGIR4mj4hz/Kt7eP2geQWqKK5yM+LuDXA1pNQKeU4M5eANpa3qJSybR2psqzDhu+a0K4OvNR9fRl70y5jBsgJtN9Xp0tc/tvrc7v+2jVg4zzr669pRhC11sizHEVeuPajUkjnIG4LMFzjfHTVolpjPp9jtVytRfgNEASBlZdZrZoSXgfCkx5ubm4QxzF+fP+BJE0ukmYErHM1HAxxe3sLxhjm8zmKsrgIt+0lQZFCctYoiAVYJ7rIi4ukvhvdoi5QhLftGELYlpFUDHlMS8RtOMkpbFR5VqXpT9MnTKdTF9oOggBhGNrFs/Jsqb3ZtRiwa4AxBqUuG6Hjc+6xqwwsFRbzhZN3AV/3uHYkZSqNry2C+0LujLFGlLCub3gJA8LZOkpIuoWXRL2ghcjfdcfwPYzrSy+8+/iH14i9536h4GE7NX3N92sbyKbUo/SmtBkM6UnnHO6zc9cWKQSwlu4ylTyNkNDQTkd3Ops2eugeAsYY7u7vMBlPkKUZvn//DlVezi4yxvDh4wd4voenxycUeWFlczo4Jo0xTpia+JthFOLm5gY3NzeukPDPL3/i4cfD0cdvb2zbhU+XGo/1oA9gM4XG2EyWJ86vizjNKaxdOGkdkVRH3QHUSgMcay5WxyZq+1x8329wLZ57fxdRd1AYZ2CGgenmee8LjyujXDsgeqZKK5jSYDQa4f7DPZRS+P79O9IkBRfNHXvbSSQdqzAI8enzJ0RRhCzLrBZkLXVE6eNz7jHt+rI0O3uX157g1AuZMYZBPACXfIPfdEwVX6fG0q7hYKzOXIPUbLSVTKlQj1oRn/Oca7vEYrIt4ngxg7xRyESv70pn1nh11Z82ZXDjO7ZpIjbO4Ti+YhfA2FoQmH6m5+SugTIfO67daFutTB2RPM9z2n5UiJEXObIsswGIjqtfEBwvtLof1OEFEvCl7VWcZZlNLR84jAUX8HwPk/EEnz9/RpZleHx8hJDCccFPPdf68/GkB600VssVfvz4gVWy6uyYdEETWB3MMAxdS8Esy1w/4cFggMVi4eR8jjn+eDzG7d2t64xC8j3DwRBhEKJUJdI0xePDml946P2icULOK/28WCzW0eYdLWePwcmcQpc2ZOs2LkVu9eLIG9dGI0szKwrJmRNE7ioYY4ijGIvlwvb5vdJqZM64m7j1iNYh2FYYIoVEEAaYjCfgnOPp6ckSjKuCk33OUJ7n1pm8u7dcxDTFYrGwky5LXaPwS8AYWwBybkXzNpCDXBa2pV7IwxdzPHps3kvj/td45XXROCV65rVXtpySLfoy6zeaC9Q3NmpQuq0Hd0kwzsCN3YSScyilhPKUK47L8/xiqdG3AtlvKSVub2/h+z6Wy2Wjy9Y+ULbo9uYWHz5+QLJKrMO2Wl3UNjLGoLTC129fwRhzmn9dHI9uo8hsoGIwGEB6Ej9+/MDj4yOUUphMJphMJrY24sh1iShXdSoAbViEELZoyJmAdRHjKc/CZWp183iUlT0XZ6/IVGUkheWKFUXRUK8nYcuuL5iMMdzd3mE0HuGf//wnkiRpaPB1bfdTr7jd+nu658/svg8BFxxRGGE0GkEp5WgC23g9bVBPUwOD5XJpOSeFraxrRyxPLjZh9n6QCPaLgNlFCcx2Y/CUZ5XkG1yyHudiazrZ/a/xyqtg22Nltf8fhUs4hIDbjF+jJh9nHBqb0ULCcxXo9QgJFWdobWlJUkq7/rxB4IFs2UVoMNVm2/MsF1AKicVycXBVdVnYDkxSWiHpP7/8idVq9SLFH9RiFIDLGJ6LbRz4dgbq6GPWNvCe52E8GkMIgflsjqfHJwCWuzkZT06iZIyGI+R5jsVi4RzvKIoAY53Qh4cHlMrSroqyOMkhrDuc9WsiXKpA5myncDabocgL5EXuSqUFF/A9H57nuZRbBzcPDnWn1fd9q33Xks/p0qLvzoVkZ4jUa9BcLCridttQHTN4GLMSMqPxCGDA0+MTklXiUoXP8faklEjTFF+/fgUDQ5ZntpKZr0v/TzVUZCg4eMP5ZWDQuLwBdM61qYkus26NjWvGzvtomv94LVOydvjX37/LF1unkbcfyX56fZxnvnj/W1obPbcQv6Nh6Gy2WVeYF0XRkOZ6K5ybOWCMIfBtWzvOOeaLuZXuOtDZpZZ2379/hzf1MF/Mt372XLultI3Qhr6VF6P7f7Y93LYRO7MAjbquAYDv+QjCAHmeI0nsWuYHvvt9mqbI8uyo42dZZnVsqwhjntn2c+TIcsGBEm7unrPm1f8GLr/+HOUUbhvseZ47x88tyEYjjGx6bTFfrNsWdUi3yIVcud1hUlWbEMIKNBfSRcPI6GqjX/RhHAsqCAHWjmGd4+VkaVqnuc9JbHP7PM/Dxw8fcXt7a/sfz2ZrQecDG36T7Ez9u3ZNikMdVoOas1tF8aIoAmMMaZKerSMIbElhVg620VbJXwrZ6Ct7zHh4a97dW+GU635dV7CGI051beif+RB7viUVA9vbn7ruBJJWIf391jZpH+ge1aNqzy2Q+66H5GrAbPVokVunxBjzqnzChl5kjRt4jC2rw5Mebu9ucX9v+dvLxRJ5nq/X0GemAukGJmmCJE0ANJ2qSxY83N7cIggDLJdLcMbd9516vH2BmLM2+8zKoXHGMZ6MEYURHh4ekOdVMKviGDLGkKXZ0cU4dcmZNEnh+R6iKEIURchzq96xWq0AYKto+KHPpB5df6m5flHFZoochVGI0WgEoNo9lOqsBtMvAcas0HYYWLKpgbEdPBjDaDRCEARQSiFZ2VZDYIApu+MQ2oBVLQTNLLmYKoS11s5xai9Cx5x7GIa4vbtFmqR4enpyFcPkcHbimVLkhK0Xyxf7quo7lLI9l6ktV5e5slcJtvGPCqaRvjUMwEU2m9ahO2XoWNog2xElBCjb676mx0VAnDYS8C/KwhHt39w+nwFyKMqixHwxx2q1shW9elPt4Vhc8r4wZlVGBoMB0iS9KJdzG7cdDOCan+QYUgAliAMMBkMYANNZRYOqqAee9JxdPwX1jQh15UlWVp6v3onmXMf8pdLGhIu38fA8D5PJBMPB0KmbtyvOugIpJW7vbjEZT6CNRhRFMNrg7vbOChUrbYW31WlCny8FisgC9pzo/kpppQsAuB0zcN4gLIoCP378QLJKMJ1OXbFQZxxCYGPXtG3SUKuoc76jDmrf6Hmeiwp05X5cPehWsxZ7r5FWrd1rKuZopXudahZjtb/tQZpzwthaEGy6oAefMmuc6fb3YHeUsPHqOxlGhygO7FsvOLNdHLzIs+3WStVYa94KZ6dlSxsdXK1WWMwXrsDkXIfwkjDGtisNwgBCCJc6Ldhxkjkbx6V0az2jVE1MxhiYYIDCSUEmA7txWCzmeHp6xHw+B0zVorfqu12q0nEkTzl3mt8kvfb49IjJZHLS8XaBsyoIsSUDKLg4235c1ilkwHA0xHg0Rpqllm94gTTeS4HzKmTMGZbTJZJV4lLhQRBgNBrZTiE7skJ1A/+Wk5UWOCFspJDS9adGr+rXlSYp/vPv/+noAapU7lqPjavUnbdtBu5UkjJjrLFLI0oAzGbK/1RsO4ZzDKX3PA/sgjgk5XaRzde2a2LN59R0uA5YEOu/3pltZZs/GlipFmbA1uIurgilTg7nTAAMUJracVFxAgOYqXhodrExbnzYSN8Z2wY8NwDYQe/C8yfR4hS6l+kCXtEfYmAwO+R4ABxAnzzdhjLOnCRaVmQuUvXaDmHdGTil+rb9HPM8x/cf3+2xayLQ9WDAc+fjjr2FAnMuyJH3pOc6afm+bzNV0nbXSNMU1LbwKBj7XBvdbszaCSWqUM0EHARaI4q8wJcvX1zLVk96zg+QnkSSJK7by1GnXVGLOOMuOJNlGfKskriD7U98qYwSjTnKDF5Se/Ky6WMwRGEEMODHjx+2w8mW6rGugLgnRWEHitIKRWFTgjeTGwwGg42iDsJGhZR5O8eQCjdIWJpS9qdGCLdWgNa5lDht9XTOJDktrXt2TIuhttQOTW4AruUiA7P9QpMUCpuCqs/dm+cMqNE2JUH33joZrzMGnouuXGyebRxm0xE5xjE09V8dcYr1QJxbfmtRQwOG0igoreH7VkqqKEtX+EZRQmMAwwwYq5xIw2DAK65W1YP7xEf43D13C/ohX9BytDY6I1RzsM4hdr/blnp7IdQdoq2/f+Zaz43ee57X2BC8Ba+yscFtbZoOxYbzpjcdu0OP237fJbsvMWadNc44hsMh4ihGqUrc3t5CCukqwP/zH/+JoiiQJMnG55+DC27ocuO5MmY3Iaekj6nTh8rUesww69AOh0PAwFVpHwtqLSt9ieFoCE96+Pb4DdKzLhYVQ12SZsSY5dELLrBcLi+iUQi8QKSwKAs8PT25qmSYaiA4p78b4W+gKfT43HltGL+O+LYuQljt0JRWLlLYRWi9bqZ+0egaw/qYFciwvtQiYWBQqhJccfjcPylK0ONwbHuKNIQ45/BbxQWRH7h/a1NVDjveaRWxhrHRQqahNUksvdQztGfbEdNx9RDcFg6oUl1sQTwVl8p6bMO5x1LKZnecU3VOerfacEpPuiwbyqrbExR830cU2wKLcztKkQYnacS6VDLgHKxTbbsQwgYOmG1G4Ae+bSOY2BaAx94jOpcoijAajpDlGbI8Q+Db9PrFUTNTQtaOf4FhdxGnsB7WXiwW0Fo32vHUI0td4hTWq3B3ahOxmlPbMWteL6zQSqM03W5EzhnHYDSAUmotan6mw+YqL8E2nGFKbdQNySVhjHH8Si30urMPNiN1XX0m14njI2F823uM9Q0NAM32FIpcDMYGAA/4omPGS8N2ddBOvRSoQrtU5cFKCC+FrmbEOOMYToZWGzbPNqTWjgXZNs/zEEYh0jTFcmn5j5xx3N3fuQxblmVn34d6pFAbDW7WG7+z1w7YFPh4MobneZhNZ8jyzBVpHuOM07mQBu9ytbQBGymcL3SynE7bkWfNTQjx2i81/i8TKazl+euNpNvefddgjHFl4m1VcD/wbSToBH7Ba6G+ELR78L6ERl+j5/Uh51d7P+eW+3MzuUFe5E5ioV7K7z5T/959g4etuSKcc6RZalX1a6/RjuqlFgxjbLSQlQxhENoJe0A17CUjCVsOfrnnv0Hva46turHb9p3n33OKrF3eqV4Hqlk1Zoxz9C89f+hopwXHW05wLXXc+A6SQ6Ec/SvY3WdtTfsc9r61dT1b3kzfR63titLK0Fx7F5M66s+1LnFzDEgv0PM9DEdDMMbwxx9/NIruSGu2nX7fB6L9hGGIMAyxXC4xfZo6vb/hcIjADxyNqS0N9Gy2jaERAdygTZDzc2ZWhvySwXDg2twtl8uTo5tU/JGlGZ6MLbAdjobwfd854+c4hrTZoyppKaXj0wIVp1PaDirLxfKse3OWU1gfSJxxxwUoSps2VlptlUTpCowx+PHjh/u305fiHHEcI89z228S3Y/0uPQALdqXopTVCkNO5RFyzq32o5DwPMv9o043bd3HY7iLlDrnYi2kXZblOkKIPRHgC4GciCIvEAZho2ND+1z3/XzpczorGtB6Jocee9vvNu59RyIoTVRFJrXxd3HH8EinZfMeNxdTpwpbn5+0R2wt8Icu+KfiqOOeeQr0jHzfR1naDhG04AL7x+41oHHOzKbIqWjwkOthzPLLlVKgQgTGGMbjMX7//XdIT8LkLR3FI28TY7aXL/Hx82K9wadKZKVUo+3b1uvbdmxYzqKCWlPPKjTSsGdSjwQXGA1t+1XBBZaLJZarpeUdnnBcxpjrnZznuStwpDUpSZKzKA7UpMH3fQwGg0YwRQqJ4XAILuz9Xy3P6z99kUih0QZMMozGI/i+j+l06kLHXZ2Y5DyR00fnqrXGIB5ACIHZbGajQB29hjpezPGuDiuEwHAwhDEGs9ns4HMiI8U5d4MWQFOct8KxBp2MnhTSpZD2FTscEok4BVprgNvUgR/4W7/vZ+UatiOFF02j1fYhL3f3mmnjOqG9Lut0/tfwqiDhUBxJpEdTOPlnBEVj6PooQnhMpOvSuDSPuD6XhBQYDAfQWlutwsrR2/v5Ku1J0mTaaFeM4/s+tNYIgsA5LYeIYdfBwDAcDhFFkZXMWSxscwJWKxAprLMuhGhWxR7waNzzMy8biPE8D3d3dxgMB1gsFniaPm1S3o5EowkE58izHEVe2PZ25emydu1zKcvSFvV40vVXLsrCyTKdi8v0PoYtFx8MBoij2LaJSddOYWejbAaunQ2RTrXRiAcxPM+zyuZKNSJP7wEUFWSWvOC6vNze3gIAlqvlwYMviiLXh1N6EmB2Qo7HY1vtlaxsE/vaAnzoxKFdkpDCtYGqcwy3vX/jOi8ErTXyIrdOocHGhqizc6DT2J2WfknUU17nSDsRnLMGHBgpNSdXQP/MYJxBK+1aZNKzadMZXtMxvMT61uavUYRJSIHBYOBapx3iGJKjNxqNEEahs9+e9PDp0ycURYEiL5CkSUND+FBwwRFGIYQUmM6mrrmDlNKlL9PUdpQSQhwdHXutuS49adPGaYZvX79tVUo5B5xx5wi6YpkzNg/1Z75YLCCEQBRGri3varlCXuTuO8/BZQpNqpSr4DZcTOlC196utvt5zTTaPjTapMEaGCEE4jjG7c2tI+ZSCX6XQXy/uoE6NXJoTK2PsrGThxZJLjg86VmehMnczn3foimEwKfPnxydQErpuCdxFGO+mOPh4cESlTk/amIaU3UxMNo1i+ecuzA+PeNLNKk/BJQqOIV/2SUc4sy2Hfh6hO2yc/ptbiKN+ctFCqv7dFC0cFvRC6v/1t5jtn658dpPgjZ9hGy053k2AlNLG7vPvNJ6YsxaPktKebKYv+OCs3WkiWwY6a36nu2axBkHRJWZ2PFVDLa44e7uDuPJGHlue/BKKXF3dwejDbIsw9dvX5Em6VFONK3zeZ7jx/cfWCUra++qrFsYhpBSYpWsXPr44PtQC0TUbSd9J3FIlVJnUzsYYyiLEl+/fUWe5ZjNZ47O5M7lTNA6Wi8GvYQpI7oEZ1ZbkdL1VOBSH5en4mynkHhdpAWmtEIYhjZErbWrTFJKOcegKyAjA8A5FJ8+fkIcx/jn7/9ElmUXbyHzEiBnkDgcdK9PBRkKIdf6e844Ce64I4dMnlKVCMMQi8UCi8UCSZKAMYblcgnStaQFWHCxtS/kzvOEaajP08JYpwKoUjUKWl4SRtvzCSoplJ8hZbzBWTPr69rmGP5MqPN2tkWkDsX6vuwZERu/2F9gZf9qOeIU3f+J0I6g0aYySZINp/A1HUL3ndxmKwpdnMZFwzqbRk4EBVikkK6FZlmUzi4/F3Xigjsay2w2s+NXaZfevbm9sevelmKlnedZswMk3VJXWpBCOs3C1Wp1VISQpGccJxZrGgRjVv7G93wUhW1jeLZTCFsZ/eXPL+s5Uzltl3II6e+LHI94NAzOCZdSwvd9l6klncRD1+V9uIxTyIVt6+J58DwPvue7BzuIB/j2/RsWiwWklDZk3VENvclkgjAK8e3bNzz8eFiHfzuey6lPTC64S3ufApd+ZQyTycSlLoIgcIZmNBwhz3MkaYJUpXuPR0Tp1XKFx8dHt2vNsgyDwQCeZ4WG2xqDB2GjhmF97oxXhSeqvMju6RBoo9eplNYu+WdzmAgXnRsdnGbbHEPaQAohLJ9qC+qpYoMDhvaWKl1aKNsRM+co/ZxDaieoe0NZlht8z7eYX3V7c+5xAPu8fd+2WzMwLrjCGMNgaLX0lFKuF/IuUHVumqb49u2bcxQEF/B8Dze3N43vPQTuXuuakwI7FpVRiOIIQRAgWSUuYnUIB3Lje2pGoN6UwcDYApYTNAR3XYsrgq0Tly+wsXqJYABtBgDr9AdB4Lic9Y0hZxzKnBd4u4hTyAV3TmFe5HZXIoVLx0Zh5CJDXQaVpX///h1Zmr316RwFiuz5vt1R1Z3CoyvAmJUy+Pz5cxWilmAMVTs3hl9/+w1FnuNp+oRv374hTXY7hsSnoEWUDAaAl4ne1Sa1Vrqx43wNaGUdQ5J7WJ9Wt8d+l3ChTMvFQLSGdqptX0UoY3BOobueIy7KwErL0ALMzGXGz7UWojBmoyOUHXjrwEIjLbgFx9hcp/0nPdzf32M4Gro1NAgChIGVf6HMx9///ncsFoudx6ONqaMTGTtWOVtLdJ0ywVzbulq2QAqbOo+jGH7gY7m0FbzkcJ0z1ihqSud/KUWAbe333BpxIcfwkmhHhgWv1vmysI5+pVN4qXXuIk6h53nwfA9FWeDx4RGrZIUoinB/f29TadVNJt5XV4xS+zwWi4WVoUnSi/ILLg3im2iloZQCN7ay101CA9cXtFTl5s5lS4St+Wv7hsV8gSIvIKVEFEcIwxCrVYLFYoGyKJCskmd37NRiidLCnHOkaWojhFW4Pk3T7dWebe9gz2QlXgulubM8c8d7zfGmjXaVd0EQuMgG8HrRDA5+8m61Pd7rKWLXprB6BkEQ4O7uDnd3d5jP5wcpDrz0bNrXhrf5xuOPXaea0N/tQoN6FK/hx+24r8+dI6v91/5eSiN9/PjR6sKVBZaLJYqicJQepRSiKHLFXK9Bo3hJqFJtrQp/zXlO9564y0SvoWpocjga57PP5pp1CrUoCuSZfVZSW1tG0UFaP5/LApFGIdlUBqvnaIzBeDJ2PLSj1QJMMyXKOYc2GoPhAJPJBFpp27xCbbn+PWikb7G2N4ClH5XKpkxfgnpG0TXCJaJ8ZBMuNh6ZpSZprd1azIWlUIRR6DR5HZ9en1f8dJFCk8APEPgB0iTFcrW0izwqTpdWjg/RJT5hG8aYRlpCsBdoTXMh0G6NCno8z3MLBAB4vgdprJHKi3zzAKz9Y423U6X9jTaYTqeOw/Px48dqccnw+PjgjBS1UNp1PKWtQcuyDKpUzlCFga1gy/PcLmJVmrkOIh+745rtRHrHreJrXa5GlPCVd31UcBKG4YY492vhmGtupGxY0/lwXEJU0QZhaQXj8RhBELh/r1arN9/s7XIId5rHI053Y+O0J9pdMaR2H77t0Oz94s03uLRyFUkZjob4WH6ENhqL+QLL5RKLpZUKCfwAaZq6Ao23jrCdDGbnVVEW3biG1sMVQtiIH2eWx2xaUa09NpegSoXZbIZVsoIQAuPx2CkrfPv6zSosVJvOfZBSYjqdArDjk4ozOLcZPaWsdInRm9HvQ50Zeo/nebi9vQXjDPP5HIvlwkUlj7FBDLancX2sG2NerH2hFHIti9Zyds/FpWWK6JjSlxjEA2dvV8kKQRi439P9Pvf7z3YKhRCIIlsssEpWGxybLMscj7C9q+4SGGMYjUYoyxJ5lnf2PAE70T3pIQhtasHzrQ4V8f9Il6ooCsstydKDr4ccLK01ssy2oovCyPZXrML4aZralPEBc74oCjw8PLi0MYlZ+76POIrx7fs39/rJuysGd0ySAqANyFukAQyMK3B5kb6XrwRy4PMsh5ACN5MbfP7LJwyHAwBwgvV1nl3nsLEYv0Zq+oBRx5r/rJ/TxjyoVWLS7+lnysAUZWHln4TE7d0tklWCx8dHPD49oigKJwtVFMWr2rZtDsep30+brS7YZrKTjlNYcT9JSL9eAHcotNEoCltVHUahKzRxG3X6e8/100bhx4NtyiCEQK5ycG55aL7vu3X6nGgWpfMHAxslzLIMDw8PNop5ofTrSxbqKa0AhXWBFlsX/Gy7v2+64a12mC5VDFuo6VL5Zl1owvj5PtbZTqHv+zaCVOTI0mzjhPI8d6m8DqXpAcCRb5W25fP/+i//itlshm/fvyFJEqeH1TUYY1xFWsYylxqII6uvmGe543TUWxkdAyrSkFJiMpkg8AMb7S2tk0CROa313p0JpUMYb6bApCctcbpcpzGONVL1dKYQwhG0qdXiW/JClLYL2LU6hfScAt+miG9ubjAajuD5ll+qtaUuUKSXnMKzdtw7PLZtT/Fks/cKXuFBDqGrtMTG/NyYr/vOudoQ0QZExtakS2l12O7u7/CPf/wDRVEgTdO3d9yPuP/1+U3pw3qP4y44h8A6MkNdJ04BRX9J89f3fUgpkWe5C6po9by8ljYaqlCNIkkKGPieD9/zMV/M7ZqB4+6jc36rzch4PMbt7S0451jMF0jSxN2PawAXHHEUI45jKK2wmC8cH3LbevZm11Wlj7M8AxZAmqZIVglGo1FDOqtesHQOznYKwzCE9Gy4Os1S572GYYg4ivH4+Lje5ehuRRO0smrvSitbNe37TpfPGMuDo/6CjLFGSuAt0pIEOjelFNLMpoYCP4AJjTP+eZ7v3Pkccu5kMMIwxHAwBADXy9Lx5CrC8r7j0bMng+d5HpRS+PTpExhjzpCcumtlsEUxQRCASOiqPL7qbeuxT6nOq0ARVTfeX3GoHHsf6wsZ7To96eHT50+4ublBHMduIyKlQFHkeHx8xNPTk0tPkSbpszhE87PB4d/FIXV1HBuf24m3diIaDpE9WQ77Gm+cvC3PaoDXnEYNMGbAjAFjBmVZ4D/+49+xWCzw22+/4vbmFoxJCMHheQL/83/+T6Rpiv/j//g/NtpAviYc16qVtmu/x8HYzRVJb5CSwFvTFDbAgCK3laD1TNmh59lYV8DgMQ+D2CozCGmVPbioKnCV2phnDU5cjfrROA8GjEYj2xt3uTw7LUu6iQwMj4+PmM/nVuvvDEO3rTClnUU6dd11epD117TloN/e3sIY44JaTLON9L9bxyq8qlQdbSCNXd/yPIfv+wijEEEYYLVcueAKjY1988qYqvhzxzWcbR1WqxW+fv3akJohkr022qYuq4XAaAPDOjSpq7Cx4AJxFCOKInz//h1lWVono4qMtbmQ9Sqlt0Ld2SLNIsaZ44k0DEeb5PycQ1gNKN/zMR6PEcexkxSq0wAOrYhsVOEyho8fPiIMQ/z48cOmuE8l5hrAMLvZIGNJUcK3htGWo0risdcEKtgZj8eYTCZug8GYXQAeHn7g6ekJq9UKo9HIpcoutmCbC0+tt3YGN2BjS81X2j81I4WNwGHr5iTJCmma4OHhB6bTJ9zd3eHz58+4u7urCg0EPn36hLIo8X/+v//P7jhWB0QNiSNMdIyuRQkJdD6n2B4G5jQKSbEjDENkeYZSlbYpRFVoQEUmu54fZ3wjmsgZRxRGuLm5QV7ktg+v2e48HHzO3BavzGYzLJYLZNnl1Tqo8l4wsS5EOfV80SyUo40JRQWpGJKybsAbp4xroGdF454kz7Isc3Q3Kig16nnjyVjF39yBiziFSZI4YUxjjI3chJbgnCTJ2gh14x47UBseLjjG4zE830MURbi9vbVp2DzHcrHEfDGHUqqzi7vn2fPmgttG4m0e1Qm7K8YYwijE3d0dwID5Yo7hcLgms+7hX+yD7/v4+OmjVdX/+nXdAeTI49S1suqdczqzWFTE+LIoHccT6I6h2QfGGEpVIlkluLu9gyoVsjzD48Mj/vzzDxTlWkXgFJL6+4Vd2S6dwV4ul64wYbWyeqDL5RIPDw/49ddfMZncIk1TfPj4Ab/Of8WXP7+AieY8fimcwylkvJKhMcYVmHRlfLnKY9S4nmd2vmJgCIMQk5sJGGOYz+aIQqv64Hhve6g6uxCGIT5//gwpJf788uc6Inbks2/MeQOX2n4pnipRUki8mpygU1GPVFNvaFLBgFn3bjbabEQKOzPuqvOgjmtAs0iGupHVbfOxz+Yybe7QnPie5yHwA6xWK1cp1ZnFugZeNannzPZtLosS9x/ucXd/Zwm6eY6vX77CGIPlavnWp7sT1HfSTdozvG8aYIEfYDgcwvd9PD4+QinlVOUJGxV2eN4B/XD/AUII/POf/2zoTh3LJax/r9JWpoIMdVc4LZTyKooC3Oedok7sRMVRy/McX75+weRmgii0wrRKKXz/8Q0G2hkd0kMDtjsYXTCmx57DS9mql6IzKrWWaaGWYADw/ft3zGYz/D/+7/9PF3H79OmTFeZXZSeejQOrPSezTnEJIVxrr65FCdub0FPPi7RcpZSIogiBHyBJE6xWK5dGJgoTF/yoaCRjDB8+fMCvv/2Kv//H320xSJX5Ovl8K4oJKU+82POoDiulRBAEKMtywymsp3WfS+nSuuBJz1Gi6mLhg8HAZcOyLDupWOjSqI95+jtJLOXKydBsK0A7Y25fxCmkNKYqFaSQGI/G4JxjuVyiKAuniXTuyV4axFeJogiTyQSPT9b5ofCsEALxIIZ4FJ06bwBOh8z3fQwHQ6SpFZAmgVfCqRM2CAPc3d4hS21VGWfc9i725DoSueXQbe5FG6vVCg8PD45LCBy/aBP3hL6rUUHWAYfQ3fOqWrssSwR+sOZSvfT3a+PSTlEcufRvWVjNrzqfiKolAbhqSnIMsyzDjx8/8K//8q/Ii8KNtR8P392miTou0Oc3eDsdWcDrOGS8HXLe59iEY/mq295PVa71Th9UdALAvfb777/jb3/7G5arJaIwwmg0wpcvXxBG4dnXcci5t//tImoMjTlRX9y01m6jmxf5Tq7Ua8Px2qpoGdmf9tp2dMEJsw7KaDQCYDViqVBwWweXfWg7R0/TJ7C/M/z48cPxnM9+5gZb5c4uwbUjR5NaqpIsGqV66Tu0bhaEbEubN37mHKPRCP/lv/4XDAYDu37Uorvj0dhpLf/55c+d3YpeG64zDEej+NVVwPOm/M9WulsL28Ys4TIdTSjixjniQQzpSSyWC1t4ok6LBr0GqPvH/d09wjDEf/z9PzCfz61C+yDGv/7LvzoldSHEya3jLg0Gyx3U0PAD3y0EjDG7oyYO5wkGlAZZnuX488ufrop3PBlDcKuZRZNxWyXcc894sbD8Ey6s+HbXxsQlQfIAWlm9ToHXqUTmgiPyI2itMZvNEASBkwQKwxCTycS91xiD5XKJ+WxuIxXDyKUlXO/yZAUpPUjpIYojyJncKw3SxbTLsXguInVqaubS53IIZWK+mENpBc4Foii0x3vpEuxDsIuXXdvgkURLF0BrHWUkLkVZoZRwmtm2dFxYRzCOY4ABSZo4nddTntvj46PlEarL9MY1xq49L0EXIYeQNjp0j7XRrisW8Svb68+z51Ldy69fvwKw4vuj0QhxHKPILT+yKAvMZ3NbONQBUB9sxizvlIpiOeNuQ69KhVJfLvJ/vlNIFUMMiGLLxxNCYDab2eKTSj8HOG2B2LbzcNVIYBUJ+/QwuOACHz58QJqlSNPUCW0LLuzkLKyT1SWnkCKzvu/D8zysEisOHUXR+j0n3hOafKUq8f3bd/i+j5vbG3y4/2A1rlarjd3/oc+VM+4cQjKml0wH1XdLb51monuitbaq/EUJKWyaH3h5Z8LNS2NloYbDIX795Vf85Ze/bMjk5HmOf/+3f8c//vkPPDw8IBoNwKQAU8AyWeHh6QmfP3+G4HZzMJ/P8PDw4DYQ7xnHOod0v96iGGpXxOCto28AXFQdqIr/pF0Ii7w4mXd8SdQdQilsNoYi7udGxxhj4LCO4Gw2g+d7GI/HuLu9QxzHeJo+rak2J6z7UtiKY9/3L7aOvQiHsOYQUjcorawSAue2WEZK6Spwj/WPi6JAURT49u0bsizDYDBwUmbL1RJfv3114406cL01XIaVM3jcc5sRsr1CCMBvfiZZJY2fn5MxauNsp5AI/3Ec4/b2FlEYYbFYYDFfuIox4LIRg3rp+jk7XqMNxuMxhqMh/vjjD5vurtJkjNuq5FKVzlHqCrS2E2U8HkNKidlsBqWU5Umc4SQDa56lJz2nLUnSI1JK23OzViJ/COqOI+Os2QbpBe18O5X9qjICFWgxo3ZN9XTtS0ErjVVuuyJMbib4X/6X/wXD4dC1GKwvCozZNpX/6//2v2Jyc4P/6//6/1h9RSnBhUBZllgs5ri7u3UcwjiOMZ1OnWPv0oJdKvT5yXHMGBrEA0ghkSQJktXbV+Zvg4FxGQgSbe6SWDUAWwlbBQvajtU5Y5+qX4UQtpew0VgtV5h6U9soIK01HzjgK2hsKK0c55e6PWmlt1YonwrqlHIpUBOCMAzdvQiCwHJiQ1sAt1qtnC07ZnNljHF8VTqm7/t281EUyFLLI6RIcFfGXZqlbr0fDocIwsDRxwA4eh7h3//t38/6vrOdQqUUYGwoNo5i5HmO+XyOvMgbvWePXQjbC3jj86wKuVcPGTjNOfQDH3/729+gtbZp4ypVWhS2OwC1jaJ2bl1JhXFu+X1/fvkTANwkKsrCkZJPBRWPpFnqOEsAbMUipZ0a8hj77wkZIFUqfPr1Ez5/+ow///wT375/c3It9WjLMfe4zSFkzGoWCiGsgHfLYFzKEB5yXm3KhFb2HmhRcaValYrn8A211m7MJkmCsizx+fNn/O1vf8P9/X2Dk0T9sKmPZuAHUFrZSsdBjP/63/4b/v6ff4fRBknVCWc+n2M+XyCOYwgpcffhHt8fHzCdThHrgev7SjvYrsyTc/GS17Fvjh66GOV5juFgCClsOj/LMlupCriK0DAM8V/+639BURYIwxDL5RJP0yeEYXjwwkcVmnlh+YtFXiDPc1fgVr9PuyKnDUpBbaw35gGDy8qQ+sNLtTk7BUYb5CqHyY3r5kPND04+JpqbqqK0aUulFL5+/eqeEUnWHGIjiY+nS43RcIS//vWv+Pr1Kx4eH5wTJ9i6E9Gh49xt4mtvN8YgDEJ8+PABs/kMy8XyZGeKRMrLsnStGUmjkpog5HlufYvycI4lwZOey1IxxnB3d4cwDC0Xt9IjNsa4dqxdQRAEYGCNjQjR2gC4Huej0cjNc6oxOAVnO4VSSJfjLooCSZI4EetLRQlpp9P4mTGn8H5qtNBoOwnT1HI5KELoeR48z7Ml8Kp80WjWJUAV31EUIU3Sszk4roijniZuOYP0vuegjbY7bGkFtoMwcGLTvu+7Ju+HHu/Zc69Xwrcq495yoitt+7a2F9FLoF5x+te//hV//etfMRqNwJhthxRFEcqyxI8fP/D777/bpvXV3IzCCP/tv/+3amfOMZlMMPhhRefdHCgVptMnCMGteHXFdyrLEh8+3OP+/h7T6dRJU/V4eTBWdfEJfNzd3WGV2F7kWZa5IqHb21v89//+351syHg0xmw6c/zvQ4tplLJ9cuM4xv/43/4HgjDAv/3bv+Hh4cF1T7rINVXVxozboiil1Ktt5J5DO+vAuF2TKPKvTZPjdkpWYsORbtncQ50gpZVbI6UnMbmZYLVaYblcNoor6D3nRMQo1S+kcG1WzwE5ZTDYSIsqpVAUhdUOPqLwpg5qrhFEgatoLoqi03aLaANZnmE6m4LNm+uH79u6giiOLrKJOv8pMjt40zRFqUrnzWutrcI5Py9yUK8sbaOu8n4KSlXiy5cvzugBa+HtwA+QrBJ7LabbBRFaa3fPF4sFyuJl5SaOrZwUXMDzPcSDGKvVyrVGE1zA93wrqVGrUD/9xNb6Ya9V6XsojDGuEb0UNRmXC5wnca7+b///9t5su5FcyRLdAHx2ThoiIjPrVHV1dT3e/v/vuHf1a1edk1WZGQqJ4uyzA/fB3EAnRQ0cJLpC2rlyRYQGpw9wwGC2be9//3f89ttv1tVGgPhP//3f/40///wT4/GYXHuaydsYg+Vqid9//x3/43/8D4RxBKkkLq6ucD+bwRgNISXKusL9bIYgihCFIaSQxE/89g1RGNkMFB+zy+/KzwDmXbFyAmsU/uu//qttDuJO1jiOkWdUQZhOp7i5uXlxQAhQoKZrkh8ZDAYUAEiF//3//G/83//7f/H7f/1+VJfmxmbfCCudwx3HXSnhbYPL2vwsXjtxsM87VRQFhC/s/JqsEuRFvt4MNIL/p7i3nBRyHZeUKU6Euq6hNAVq3IjDSg5VVa1VJ/Y5pq5tR/fF6AKBT/OW4zg2iD/kuK+JjeSMAbI0eyAFx3N6mqYnKeWfpHzM5SmgJTtg1nZGxy4UPDHZ9LlcS2C05Un2RVVV+P79OxzloNfrWXcN3/PtJNrWx+oihKBO5OWSOJxlVcJzvQc7n2N2safgV7DrihSUjWK7O85u2Jd9j8/hHRSPgbaw9q5rODe01iirkrxNXe9kgSvfy5ubG4xGIwghEAYhkiTB//v//b+Yz+bWoYQ17QDYMXJ3d4coivDN+RUQQK/fR6/fw914DNdxoCuNLE2xWC4QhQFc10XViAlnWYrVamWz0124zz87+B5zhni1WtmMe13XVnzfcZyGQ2rg+R7+8z//k4SunT2yImItcRHHsZUgmk6nlgJyqmcupLDUirLshjPRY2hnmI7JMr1EjHrf+8u8Qa56aaMRhiGcrw5gSOw8yzNkaUZ+0q21YZfVXBusqchzl+M6tkohxUPNPG30wVxua6UnBKBhkweHJml4vQjCAIPhAFJJJEmC0WiEqqw6k5XeBc5UK6keyK75HrmvVRXJkB373pxEkoZLDLu+x9i3RMgPyFHOuutVN92qlbEpUyPJhPzQXSVnTfI8p12wUhhdjAABW2br6kLHHAz+O5e922A+ShtP6TkxB3D72dmuyXqTWPygrLLF8+PvOY5Ddk0wuLi4wGg4QpZlCIIAf33/C7e3t/sFhC19MM5eaK3tJCKFhOu4dqd1DO/nJXgJz4dfXAAb+n7HdmHzscfjMcbjMS4vLzGdThH3YroPrktNLvVa7LS9eQNo/AsBFEWJoioReD4cKcmTt5GGSFYJimEBz3VQaw0D+vkfP36Qo04zLp5cVDqa+Xlt7MuV3e7w3/4+6xNOp1Pig0ahLSkzbYA3X2m6xD/+8Q+yqnSdvZ4Bc9CuLq9weXFpm9Am08bvdmvDfMxcyYHsfD7foJV0EZ7nnUwTtc0VbGeGuMOUN/7Wpm1rjt1GHMd2LMRxjCiMEMcxAJq/i6LAfD7HH3/+AZ1vrgW7KDcbGnh1bY9nP6MX2+ceRRG0IbtRK211QEJCOQqD/gCe79kqHh/nsWzYU8fm9SIMQ1xeXsJRjk36wKyP3e6B6ILmLbB+p7gi4PmbdfUwIC3aOIqt8w/jEGrdqzmjnzqQ4ih/I50qsPEA970B24OIOFLX6Pf7yPMcaZZ2ere6Dw7l1vH91lpbseyNDYDAk6UTntSiKAJA4tUwsNyh7c96MekZxOdxlGPFxttlsTAMyZ+zLEnjqzivnJAljDclkLqqT1ZuYSN6IcmbeDgckjJ/rfH121f81+//RRzfHbqQQgh4roc0y1CWFTzfQ1FtlQOb96woi0YA2YejHJSmxGQ6ha5r/PLLL9YN4BOvC36nwjBEnueYL+ZQDnnmctNPlmXI8xyr1QqTyQx1XVsy/T50GyEEPM/D5dWlFbtO09R6xJ+y85RpMG1/3y4Hhq8BzvC1N9vbTY7PBSt836IospJlZVlS4sBzH6x7+6wNnku0hMFgYJvVeB7vD/qWK75cLvHnX38eFAdIKW2GM89zm0wgoZNN+7aXrvl2wwSqBM7nc9xP7uk4MBtWpF3CdnKmrEoMR8ON5A/Ts4IwQDHfbLA8KFF23Cm/HYQQDyJgdl8wouEu6uMmkTAIcX11Ddd18deff3V+t/oW4N1qr9dDEAS2S9vCPD2RMBG73+/DwODm5gZ5lpNw6KCPKIwOPjfOgmqjIYyAqdcZzbquAY0N8fRzox0YWicKJqofGkyZzaz6bDpDskqoVKxrXF9fk61Zo70lzUNJHM4EU0Zi6zwEuTNooVGVFRbzBXpRjCiKSJDbUUhWKyyXSwyHQ+tD/dHwkkzxqVDX5MTk+z6WyyWShJ43P8MkSfD9+3dL7VGKGruMMUiSxPq+vgTGGPR6PQwHQ1tFmEwnmM/nBytLtNH+Xa1pjLFWbFcrNK8JlqYREPYZs1Taxs+1AqIHSh1No06v14Pne/j9998xn88hpcTl5SW+XH/Z/Pl9stjNRjvNUqJ1aQ3HJY50VVXIixy1rkmjuDF92AsNL9zzKEOYl7RWbDh57BEgWxh6b4xjML4fQ9c01i4vL0n7MC/ssbuUJQRg3cTKskSWZhiPxxubMSEEojCC67gbMj2HNuCePChsZ+xO0lVqsKFrx5OFfRGOOHTbEkophS9fviAMQ8xnc9u+31VY+5+mXNq+x+3AqKxK6GoPLaftUrAgbbqL0QX6/T7SJEUlqo1n+9yCx5I5VVltGHkP5XDjGeybwdS1XjvOSJJY8AOaQLJ8LUTeJfD9Yh7usY1Y7fGvpEJRFrgb36E/ILssx3FwdX2F+Xxuf65tGcY8tF4cw3EUikbJn51xjDQQzcdIIZBnOZLVCoEfAIasofIkw2w2RxiGzY4b0LoGIECX1r6+bj2P9wYeK2EYoq5r61TTrqCwT7XWupEpym0g6Hneo8fehjGk5/bl+gt830eWk8bl7e2t5a2d6pqEIN54Ua4b+w6p/rwW2vx1YlRsWosx165dWXkxbOFL2IY75VBZdjQaAYANwi3to3Vftu8RZ/B6vR5giBrCjWf1sLa/81jg/VRApLXGcrVEkpIOahRGGI6GUEphtVxhvpjbaghXbjayXU88T05AMI2AG1cdx9lozjsYhipVRUnC1/1+n9ydDLBKDpfSeW3ws2LpsXqxzqQD1JV8fX2N/qBPndv8ewdez8mDQqUUkZNbLePHPEzOqmwEhJJS7NaUWzdt9nveAz4ODDAYDHB1dWXlaTYEQzsGIYS16PE8jwRVWzsHJpInSYLJZLKXRM1GKaHVuMHlWT/w19ZTz5SO+Rhfrr/AdV2bsVKNKDKL1PIurR0gvvRceSKuavIXtqUGYKNL61XoDAd+n8+Xm06YB3boeGPBcS4Rje/G+O233xBHMfIix+XlJf7x939Ybk7duAxVFWWcLq4u0RsMUFU1udkUJZZNRtgxioJCIYBm4V4uVgj8kMaecOB6PmazGcbjCb5+/QrX8WymgILe9f3/WbM/+z67l96H7eNKKRH4AYwxmEwmVmYkz3Pq2FTK0im0pvmRg0QuH+/zmVEYodfvQTmU1b6/vycBe/G01uJ2w8H2v9t/Z2eGdhMU8Hym403HkgGEog2y65IWKleqAGxYoabpAbSjRv+PF39e5zhIYl6w3ei2Ln17jBhj8E+//ROGwyH5HacZZZvq2mbcyrLc3QfwTKMJc/eVpOvnLJ7v+1COsvqYwO7n89R7woE3N67keY6iLBCBVBEeO+ZLwesY9yaUVYm78R0AYLFYdMbr+AEMZU9dRSVjy61s/LWDIKCssOchSZPmVw6PXU4eFLqeayUqTn2TeUDwroGDQetBueeNKMrCZrF+/fVXuJ6Lu7s7LJYLWkA7un61d4wcELRf8Lqu4XqutQfaJ+DgEhFPSI7jWNkLbWjic1zHTgDtnckuDIdDXFxcoCgK3N/fU4ahCYSCkEQ2eSLZKyhsypoc1G+YvO+41K6Vo3jXx2bvR0Fs7u7rusbd7R2cX9e762/fSDScJhQmhYe4vv6C6+truxgZY+g5aU28la3AXwjabCRJYuWE4jhGmqSWa3Z1eYUwCm1zmKV4iBfsIj6xgfaYVZIa4WpdYzqdYjwe20Cq3b1vXSy2xvtLuyulkJZndXl5SYLVTRAxm84sReDY0nEbRhsrSLwrgDw3tNFER2myYNvzCfvTckBelftpxfK9DPwAylEk8eI4YO1Gz/cgS4myKJ/t6O31eri6ukJd15hMJnR8KeA5HvzAh4FBmpAXMmc41yfysnOVSsLzPcvFK4riaH1cow1qrMdyXVFTi+d6D8T+jx0bxhgUeYFJMbGxQ5dKxm08F9e4ros4ilHkBXH2cdz9OXlQ6Ps+BoOBlRTYO5X+CLiUwEbQwFrV+5CAkJFnOQb9AYQQuPl+g7vxnVXr74r/4TZICoQcR1bL1YNr930fF6MLIhW/oCO0DX5eURRh0B8gDEN4voc4iiEkqcDHcQytNe7H91iWyyePzbIYk+nEcjQ50xmGZIlYFAWMNva5vgTse827S25caXdbdykI3EZbc4uzsKeCkALj+zEGwwHiOEZdE7dwNie+4XBI9oij0Qi9Xq8p9RAnaDqdYjqlhYSkbqqNqVJrA61rJElCDieSMlNRTILXLOt0eXFJotmNCDFbJkJ0Z6F/L+AAjDuHZ7MZptOp3XTbObD5nzd0/L/Wj5cJd82bQtKG2/M89Po9+47NZ3PiYzUCwPz+HboAtYO/ShPntWubN2Cz2Y4rYLvWtADBQZs8IZrnIIC4F6Pf70MphTCgbPxwNESvT5Jpd3d3G+Lz/Ptt8CZ7tVqRfmjT2McJEJalWb+TrXN5QWDEbi6+R/7EvEk4NijURsNUxlIipJQIQrqneZGflM7FSQTrxNSsHdsb7PcAtrsdj8cn2UidRJKm/adSJJjJNkV8kixmzRPJIeDB6DrUmVSa8qiAkLkXq2SFv77/hcVigTRNIYR4IO3SJQhB2TG2oGORcAbv9B+7z88Nes4QDkdDRGG0bh7Q2JhY0iR9wMXYPvZsNkNRFBsEWCmllTBJkuSBxuVLYYwhwVtXWX2zGo9nLrfP7dx8JSbWO8qBcI8oi0DAtIIt5vfcj++pIaSmTuerqyvSI/z1V5uZ4GebZTkmkyl+/PgBoOGe7QokBCAE+Y4mSUJd3hCI49guQuPxGGVZYjS6QL/Xo+BS181nve0939VtzdhQMtjxs695Hk/Bdvu3Ouq5o3ixWFhdwnbj0vZnOI5jRc1NQ7PxPM8GkFb/rbn89rvAMjSDwcBmabTQ5FqTrF1rBMTRiV/mAm+XM7uUJWzfJw6Id52fMZs0pg1+9nMdw6BycRRGuBhdbCRUPNeDG9N6xHaGeZ4/eqw8z/HnX39ubBaEoeYNdili7ubORsEngkQhhNU/9DyP7NQENWme6pnxxrKuayyXS2RpRg0s1WHrxC5ora3dpzEGQrcaTN5BYGgMJVH8gBJAVVVhsVzsrS6wC0cFhcx74NQ5BKzwKPNEWC7D8iCO4dQ3u2XHcawv5jELO5cr05RKX+1dKg/MTsIAla5oUDQE8vYgdl0X7JW4a3f11HUJSS4YvCPOcuJYtn93MBjQgtFoRW7sELdeKDZ0b/++53lWLHy5XNpd8naJ4Dnw4sVi3VmeQeJx3tSurttzgrmFVU3P8uBs4dY9F0LYEuMvv/xig7/RaISLiwuY5kdZrmcymSBNE2RZZkuPxhigJg1Qg5bOmFTQukZVkj+p67oIA5L/6fV6pGWYF6Sft1jg27dviCIqAdGc8PabrfbGdWMMmNbC3fr7a4yLfYNCnti11lZaht2AdnV4tzloxphGnzBtONd0HJYRKQryjuWgkT6U/zBWi+76+tp6xS6XSyyWC3pPQZvQl8y9T841gjRGi7xAWZR2Hjn3e7kLbU6b5Wa2g6cmkcA+1NvJiueePx9XKQqSp7Mp0jQFQIFzv9/HYDgAa9M+l6Edj8f272znxpJFP3782ND1fdAI0j7s1tzCCQPXdeH5Hu7H93A9Kl+eqtrRfk85SfMaQRpXHTeC444GhNubWQEBz/fw9ctXMtqYTSkeOsGm+6ig0JimxBD37Nc8jxZoLi1pQ0FXuaJSxzEdZTzp5UWOPCNi9T4lx58GgjIBcRyT9dSOtn8p5Yah/KEDva5ot2aPKygIi6KIeH0HdCCGYdjYb+X2pQew9w5HSklNNQIbPCc72XXw5d4GZwu3ievHwnVdlGWJ27tbXF5e2gnbGINVkqAoSqxWK6RpiuVyCSkFpFTwPGcHF5hPqtWxKCgj0ev1oI1GtqTgn99Hzv58//7dEuUDP4Djnv99bXfV83gxupE3eiVrtZcumO1SZVmWtqmL/9+1yePN7QavFth4VmEY2oavPM9xc3ODoiyIl9tahDlDORwNbYOK0SSMnmXZXhZ5LwErJJzE5vIVobWmbJ5DgQRviNvfl5ICjLIqD09WNHPZqpF54gBQKom4Fz9ZAXoKvudj0KdNAYuOM7af53OBPGcc2QL2Jb/3Epzr2Z9y3n0LcDW23+sj7sVYLBaYzWYot/VlD8TR5WPf9zEcDe2/ecfqeZ5Vfdc1efIe+9C1WYubMufgNWULuiSJ0AZ3Ubku6Y9tT9R8X8qyRFVXNiV+CLYV7vk4VVUhz/K9ByJzZRzHwe3ilkoCTZZwb/HxJksNwPKR7Hm/UtfxKcGLf1VXcGoiqPP1HLvwsojx/f09RqPRxgL2/ft32+BDgSBl7+r6IS9oM8gA0GSJpJCoSuIgsu9mURa0cVOSTOs1BRRVWWGplw0p/W1FxPk+bo+NbYpI++fOHRTaklYrWNvmDG40OTRdr1VVwXGcB2Ofg3LXdakBzXVxe3druWz2s5pycBAEuBhd2FLUcrXEbDZbW42eaE5kTnhbqaKr0LUGBKCg7AbuQROQVKQqcECD5UZmsTmsHQcQ9u/7WoECNFdffLlAFEdYLBZUuTGH80F5LC+XS5t04GvoKtoVAUaX14anwLqhcS9GURTWXQh4WSLEGLNZJdnC0UFhkReYTWd2kvV9H0YZpEVKMgkVtejbVO0RZFGjiZC8wYk5EQQENPRaDuDExz8l+LySJEFVVhtad8YYDAdDBGGAqiaSvzb6QXnxURjYxYW7Y3lSYvFP5RBd4CX+pMwNUQ6VRfr9PkajEbI0I+08ccRCLMiXVRd0biwV8VjZvEtoPwP2gOYA/xTWirw5467vb9++2eP6vo/pdEplpbpe82kE9w/syDY1xzRaNywQYbsYOVBQUtnnCbEZCElBgaLB6XhB+xxj14ZhWz5ju7x8yszVvsfZPq9dx2n/vSxL3N/fW49r5iNWVQXXJYqJNuuOd84AKqUst0pKcgjq9XsIwsDywBfzhaWAHPvceAyyQHNSJAfplL41hBSWBrVrfgn8gDZDRW3n5JeCm+OkoXefy+nG0IaKqSUCDQfY6J0B3QM+XPNHGIa4urwCDDaaVA55lkZT125VViiKAkEQkEQSjm8o5fdNSmmDzXajpFIkN7avIQEH3O2NnxAk8RLHMRzHwWKxOLpR5q3AcVZVVrgb35EsVatfo00JeZDUAX/LPMqNPToozPLMduvGcQzXc6GgkKYpkiSx+lkQOMlCvUtH6VRlQikkKl1Zrsspj31SmPXLWeTFmgvR7PbDMKRJvcUx2Iv0LCgInE6nlO1tZF+4bV9JZcttu2RkNoRVW13FYRji6uoKrkfeqUyWNvqwoJB3zvxx0m/cQRpR604+ux3gheZUQch2puju9g4XFxc2i/T161fc3Y0b67t6cxHZegzbi48QwjYQc1mLsxl2B2pabkMPSlNr5YD2ub4mtj+jnXVrByT8f7vU/lRQ9prYFZxu/9/+ubqusVgs7Gat3bxVFIUNKMIwhBQSF6ML6kBtPME5UHQcBxcXFxDNpriqSObCPuMDy5d8LsCaBmT0WsS9y1kmAGuKjsFOuRnfIy9z68ay59zDG+/lcmmz7paz32hPcjb4yXtlAKHWDROu6+Lb128IggDzxZwyvk2GFjhss9JucmFHpjRNN7KGh4BL09y8BmxuLFmOKcsyq1hxyLhp00cGwwECn6TR3sM4BNZWsbxGM8fVemO35vNdlRL+96tlCmFoF6Uc0lLa29amQxBCIAxCAOvU/XsALwCsH8jaUVVdWXmJl4IFvVmehHdoAOlDhmEI13PJMaQhqj81sWijEbohDAy+ffuGwXCA2Wxm6QRHWfJs/YrtWtP1uwkIGcYYm4059TuUZRmmE2o6KcsSruvhy5dr22m8Pok9D9wEkTufP39pa53gj9j1O6/xvrWz0DzW2mXLNrgsy38+N7ZfG9vB6K4Adfv8uCmEv+95HsqyRlVXmM/m6MU9SCnRH/TxtfyK29tb+x73ej1cXl5iMBgCxkAbg9l8hjRL4ShnHUwfUT4WQlj1iDRL381CDDy9mRaSNqNVXdmM1h4HpudoYAN7DiyVQ8LQzOF7indtg4LWmBiNRri8vESWZfjx4wcdH+LFmpVPnrYQVCnUFGhydvOY4zmKkkuBH+x891g/dTab2eD8uc8UUkAYsW6SagWF9n/XgSrVu8gWMvVHSbVZAXxqfG5tMp/CyXQKWQfJUY4lDb82He/BxR3ZOSSlxK+//YqqqnDz/ebhZ3W0M4l3+y5IsNpRjuVySSFhxMt3VKwVpbW2fD/uqlOOgh/4cB0Xy8WSyiTPLJqcSRxdjHB5cYmqqjCZrDULD93tbcPArDvG38caswHegUspEUXRSRdKbUhO5Ou3r5RB1QJfv37F/f09siyHlIdlf/hdeHIBXPeobH65RXdof+3Q634syGx/nSd8Dgrb3D3+ertp4zFZql3n/prYlR18KmDdPr84jq3G3XA4tDqjF6MLhAFphQZhgF7cQxRHkEJAG4MkWeHHjx8oisIKlT/oTt3zOgAyOGBZlfcSEG5jW+xYScpi1Y0rEM/JLwFvUFzXhampasBdvo7jWIk3rrq95F012sDzPVxdXQEAJpOJtbo8Zbm+qiqStzlBFZCbqzizvYvOEQQBooi4ke31+KlxZMvq/N7IzaCQEymlW3Z+k8L3paoqGGk2qhovPgbfh0dimeODQkEpZHa9yPJ1h1pZPc852+ujGu7SdhavXUPf/vnHYNOqDReK0/T9Xp+6NtWtTdHazrhtzkZH4DrN4iUAz/cAQV6OZbnu6tvgVG3dqPZ9amtbtTu7hSDOaByT9EBZ7u6w225qYekGoykT9tf3v0hwu1W6e+k9ffJnLI+4u8r0z4E7kVnQ+lTwfR+rZIX7+3tcXlyibnbLcdyzWpdP4SFdg8AB1UsmpPUxnp7ET7FQtc+prffGE/5Tgeh2BzuwziCyHeE+u+5Dzr39J/9919d3/bsNO8c14tVVVeHm5ga//varXRQ9j5QEPN+z113VFdIkxc2PG8sHtw4mR75bHGgXxWkCibOhRdR3PRdCio1r2ncc8703MHbO1IY83YejIVzHxXw+f3zta6Eoig39x+ViifvJ/bqp7wgKQBv8XtkE0JGHNMagKAvMZrO1K0878HaU7Xy2ZeUdlJddx+XYwXFIr5V92oMggJIKX79+tTJbs/mMqBUtt65zVgw20KyV7GT23Px7yAb26KBQSgnfW6e3q6oi4VuDV4m6rRJ5VT8g3PKDb+PRSazJgLHHse/41gFEKtqlsX8rw3KmhDnJBHkq8IIVhiEG/QGMJjV7JpBv47l7tLEgNQPQ9SggdF0Xq9UKedHwAZ/J1vLzWSwXMDCYTWe7CdJHojMv7YHge8Ldi6cMCrnhYDqdotfrISvI3nE0GiFJVqiesSp8Di/q0n8kY3hKbDeTsJNKe6Oz89R2BFzMV2WKQ5vwzv9vl6WfwkvH51McxscCw21sc0o5Q6qUwnK5xD/+8Q/0+32bNQzd0DYBFkWB5XKJ6WSKJE3guu7exP6nrs1RjuVCv2fwvVVKIQgCq89rv//COY0DNNYnBDZpDGEUIgxCZDmJxT8lns3guaMoCtze3lJWNsup6eDE4vHbY+1YagFAzat5nlOyppWYiFVseXL7jkdeuwVIaD+OYpQVST6VKCEFJbaCIEBRFtS88dJY4g2xTd/YiH123JNDFFRO4mgShAGkkFitVuSx6HmvloJl2Y4CBYry8IlFCiI6K6msxAZ3yda6tkryrF3GE+MDgdsuZA4FZYNGoxH8wMdsOrMOIkc3LwjaoYVBiP6gTzInk3tkaWbV+7eDSEa7gaKqGqmG7mbmzw4hqFObeH/uwYHhrndPKWr+WiwWiPu9ZsftYD6fYzKZHFY+Zu4TBys7JqCHk9Xm52xLtTw3bzz2/XbzCGcwePxv87CeK7vuOvb2BredNWwv6C895mPYh8d46DPjzW6apAjD0Fqz1bpGkRdYrpbI85xszISEbhND93x/tzMVQgpqTjxi7u4CuMGC+X6sKQmcIHssYP2Oh8MhpJKYj+dWzFqbx+d1IdZZpLomAXug+xx5gRaXt1mPubzLIGpD4//caqJk8Wng5e9ElmX466+/1p8vBYaDIQaDwVE0li5g19jY3vDuKs8zjg4KuTOqKCi6D4KAPvg1Vn+x5i7WugaO0Go0hlLJX75+ISuwigJCJcnT8Z//+Z+hpMJsPsNsOkOhiw0+zVlLyVsf6Xu+9cecz+eYL+YH6Vnt/KimzMSuFOPxGIv5ArWurXD1Y/eAd6a8UNd1vRZp/sQD2GxhddpsodbaUgym0yn6wyFmsxkWiwWSJDlNybZ5H7YnpMdKHId85nNlkrZE0naQeCzawSUHnRwYbusGbp/XPngsG3iK+8fH4XuV5zmWq6XdaLN/ba1rwAB5kVvdzEOx3QlZFuXRDQldgJLKuvmwheOpsnBCUINJHFHDRZIkmC/mVuXjqXtnjEFWrJ2JHOWgKIvO32/OmLqeizAM7XrTHucss5Rl2YYu7UY5/Yn1mJ2zAOLhJ2livyelRBiEViS+6/erje3KxXMUKiE2bVG3cZKgsKoqakk3xL9jSQQuPR4KA7PRJSUN7YCsaLU2EOplJZVdGAwHGI1GRMQuSvi+b7kzo+EIruuiqkldviiLjZfe6vycIfXV3n0PB0NcXF7A93wsFgvrPLAttbHPsbcX9rquMZvNMF/MSRuxbgj70BvnYj9vx4Bsn8fGMz1yfJzr5d13vD3HA2rDLs5NEP3c8Z49N0OToBAkHfH73/+Oqq5RVxVqrSHFHlsbsckZ3UgiGZKi2dXZuD4nJkY3J2baB9v+N2ApqkKAD0F/rrOqVVmi1howW2+jEQAEZDtIRXusbt9D+jm58/mYhs9MJ6/rGpWoAdB5OY4LpSSUcuj8Wue7Hza5l0Lw+a7/veZlPvzaxpG2nuv2uLBC6dqgNmtDgI3s7Y6N74tHS4vvJYUEJAWa+zgXPfeunIs2EkYhfN9HWZZI03RtbbfnfPTYZqqqKkxnU5RViaqsbBPddrl2FzhzzWLaz/38U9guV74meO3g91pJtTH/1ZoczKqqspW7x6gWj4FjBwAPqGHaaFsZ5K+10b4P50psGGOgQRtSR1Hgz+cshLANTsd0lx8vXs3kWgP4gY8wCK3G37H8gm0eD/MXHbX2XgSagXuAI8ZquUJVVVQ6qWr89ttvCKOQBH/H9yiKAlmekS6TWQdML3kx3wq8w0qzFNPpFFma2QDgkDT4dglQgLS35sV8Z3nwueO/6j16P5u5vWAMCbRyd/e+JdZtCLk5bpMk2fz+MSf7AqL3w18A1sz07dLy1sE4Od9k9iGwtn8rK5sx4AVid8AiNv62HsM7AimI3V9vBVi7Fn/dCEE7DgVWjuvsPM7+WN+vxzmFj2Qpn8kWvORrh2KbY8Zd3dz8dsrPOBe4MSHPc1idzhOA520+NgcyUshmV/P07/N80S6rdhVcxmRUdYU6IzH/pdx0QbsYXVAXvK43sn7tYz0FpoilWfrgZ7nRlKsAXQXfDykl4jhGr9fD+H5Mah4nethHB4XcQu65HkIRQggKItocnENKrMYYSJA8hz1Zx4EfkDp/gMCq8fM57HtPtNFW04t5IT3ZQ1mWGI/HWCUr25l8ylLUsWBOAED+s9MJ7SiZc7Lv7unJz0Kz2AkqW7Rt7Y7mK35iJ/g+K6WgHLW30fw5s6ecLWQwH217I2U3LO1Le+a0uWkkL/IHnZ777NxfY5ff5i8qRc4u20T5F51bayO8kX3fM9u/3ez11mg3TXCcXRSFFXd+zxBSWEFvzhCeeky5jkvc+aZCtY9Dyjba2fvt8zxntWX784Ve6zPWqB9kKUejEbRpvOKl2jvjLKRAWZSYzWYPYhKW/mH1hy6PUasb7DoYXYwsb5Rx7Lp8Mp3Cqq6QF6Q9VevaPrBjOHdM5GU4joPAD2xgopSypNNDUOQFyqpEEATUkRTHtizMcg1tSZquwJj1LoktkViwuU00PtXOwfM8XIwukKYpJtPJSY75iafBAQbrnu0bGL4HPMhkP5N1ZN4ydxJ2jZtqm1wM+eQ6yoHU8sXB4S5y+CHzztkb39oQdB261nZteO8wmmxcWU+QNwEnO74hK9Fe0IPWGqvV6iA/5feE7YQLr2Ntvq7V362rhsyxX0ArhEBZl1gtVw/eNUc51tr1FDajp0Y7sFdKrWkL7KBzwvM9KijcLmdwpqrNtdsOTPaZyPmFyPMcQgjrU6hrTcbeaWY/Qwq5dxBUViXCgNw2RqMR1eQrCgBZXmebzNqVwdImlfJlm/VfjgoI28+IG00GgwGCMMAqWVll/Uc7QXd0oDLiOMa///u/4/v377j9cXvwOXYdpxgntSYnCqUf6uN1BeIJjiEASLT0xLDmuvAiUBQFlFKUGWl2wPy9qq5sibiua2tfeNS5vhGqsrI6Z0KSi4fjbnZTts9pV2mYOzJ5g/fcHPQWGcJDGmeMMQ/kvd4zjDG26YGxzeHaZ53bLqEyp3gwHAAgHibbsPmBT/P7Hk0tjuPg3/7t31CWJf7+978/aMzYaAw7U+Zwm5vOVQQhBGCAKIo2nLTapgf8p8bjz4ApOUKInUGf53vwPA+z2czGG12Zb40xkI6Ersi6NfADanIKQ3genbeBgQoUxvfjB3PMvjhZphDYLFudIojiMlqtyZNTSGF3CCxGe8zxPY8kZ6IwQhzFSFOSaBBSPMgOdmWAPIdTv9Ds7FDXNWkfMgezrkmfq1nYXwohSLLoZ8x8nRLMbamrGtrR79o+8jEIQbaSrA3K3alVTQFVXdckD3VkMHgu2EWrNsjr3DpesMSTDajNejHe+f6+kLfZqQxhAy6xllVppVQ+8TRcx0UcxVYrV4AqZty8ydnXfe4lW5++N3C1cDAg/d0szVBXtW2g2QftMr8xVJKXUlq/5aKkHoKuzTVlWUKApK8GgwF++fUXKwJvYPDbP/1GLjBCwHEdjMfjoz7vpEHhqWEMCYLyzsxGwC8g274EQpBLx/X1NaSUmC/mVtn/WHPvnwVSSvi+b4NinpxgYLOq7yVgPgYPdtSv3JXHk36tKTBysdty7b3ClocUked1rVFWJZIkoUC4LS2D5xpJ3geYr+TUDtlGNtkmzoZsj7FtvPQ9s1nHhod2asHifcFZ064ttl2FkAKeT84dVVVR01LTYJVl2bPjZNfxNv6+7Ufe0WCRzyvuxYh7sW28OYn+bgPXcXExusBoSNw8NrPo0j1RUkEbDUc66PV7AGCzngZUUZFSIo5iVGX18weFVb3uwGxnl07x0LTWGA6H+PbtG+7Gd0hWCcwl7SbeM/eFF5mDgxbR+MAKIomzaj8EMBwM4bgOtNa4ubnBZDLZO0Dv0gvXZXC28L0upi95ziy9wx3FWZY9cUCclLt1FhgKkhbLhZXccFziSv8MEHK9oWb5EM4S/izgzcm2ZNqh2KAGNGoPbHUZhRHcry6kImvR+WyO6XR6Go4hUzo6Mr9wkwnLrMBQNa8X96xNalVXlHHWrfLyIZ8FA2EoC8le80maWPefLiEIgjVNzNB94rVXOQpFUSCOY/z2628nGY9HBYVPlYhPlT0yjRQF18+LvKBS0wmyNK7j4m9/+xsWywVub2+RZim1dhsDz/PeBbnXajs1LixKqXWJ4cAVlLmVNWrytJYKWZaRfaGgXYoUEr24h9VyhSzPNn63/bmj0QiD4QC+56MoClxdXUFA4F/+5V8QxzE8z8OPHz/sRHesWO6p8dyu/KU0iX3eh3anu9XiqyorSPue0O56FEJAibVjUFZklEVq/m306bs4gR0NHEd0cp4KuiaXpLIsIXLqinQ9F577kFrR1rJ7CezPnWGtl0KiMsTFdlwHVVmdzCava+DNN4/tQxbkdkDIDYRxFGM4HAIgX+UojmxTS+AHyLKMmi2fuKX/63/9L5thYncQ13Xx7//+75bj+fe//717tBRB76fvULB2dXWFfr+P+XyOLM1Q5MRn5xL6oVBSwfd9+AFVwW5ubrBYLGzQ1SUkaWI5yQCs+5DrutBGI/ADciDyfZSr42OWTmcKmU/Q6/Xge/66pHuiB+e6LlbLFSbTCVarFTzXs8EUC5N2HZxGD4PQdiWdYrcj5NrJJIoiJCmp6rP932AwgOd5FKjkj/srXl5eYjgcWg6E65H0j5QSX66/QDkO0iTFYr5AXh/voPBmeCHP6xSoa9Ltsp2O7wRSSTiSphgO+sqK5KO4Y94Ys0Ea/4gwxiAvcpLXKkrbkNJ2/+GN1jnE8l8KDoyklHaObjtP/GwQUiAKyA2rLdV1CHgTKCX5zHMCZD6fQxsN3/cxHAxfdC8vLy8xGo5sEwILX1d1hb7Th+M4mE6m8D0feZE/OOa5Np4cXAsIDIdDXF8RrWsymWA8HiNNUjuejuWk17q2Rgyr1YokhvRpMr+nhlLK2iqyHzvQ6LVWa0tU5Sjb3HYMOh8UhmGIKIygjUaWZiRRc6IxO51NIaVEURYIgxCXl5dwlIMkTWhn9og7QxcRRRGiOMJ0Mj06KDSNEG8QBLbxZrFYIFmR6HEcx0T8bconT3G9bm5u8OPHDyiHjve3v/0NUkr89ddfWCwWqOsay+WStC5f0TP7FNjQjuPr3SODc8jnAbCiv57nvaug0GhDJcS6IjmSqqY/63ovjbEPgYajq2uNqq6oG9shHjVrpR5NC3llaK0t3QSg66mrunOSXqdArWsoodDv9ylYqaqDnot112gyetz0AACr1QrL5RJlVdrNeZ7nz65JSZLg7//4O7Isg+/5uLy6xC+//II8yfH777/b5h8O4Lv4LnKVZL4gb3buvj4Vl5CD8Dxfa552tQrD/GPeVKdJSvejManQtUYQBHCUc/TmBHgHQSG7GKRJijzLN3QLj4XneVgl9OL14h7+57/9T1QlWfalado5HbSn4Ac++v2+1WDil8fqprXw3HUxh9NzPTgudcBlaYaypF0J79LyLEdZPD0Ii6IgWRUm1UNYvanZbAatNYqcOqeE020jclvWbU3+b3W+dV2jLMpOaRbuLJ23MqjcmZ4XOfKMNEw/8TR4MTTGQNbS0gZcl8SMdy1cbXmqczbicDbKcRwICGRV1un3+RgYTTIhYUAOWO1xf8i6wXMua+Yyx22VrGwGDQbIUpJk2eUuxUgSSmrw2PFcyjrmGQVA3EzBDimH6mGeGhwYCwjMZ3M7Z2R5BtdxTxa0CSEg0TS5NZt69v7uYhKI6S7aUHJgOpsiTVIIIRCERCdwHdeKcx+LTgeFAL18SZIgy8jkW2tN9XXHQZ4dt8hwB08URjAw+D//5/9Y/o7ruiQc/MIX/LW7Ubc/y+o6aQPpShLfVA6Uo+B6LvI8h6Mc8kWsNgf6S4JEbtWPogj39/eWa8mdcUIIa63TPt521tCgsf1SDoIggJBk9l5rkrRZLVe2tNwVwnMbj+l2veYkuq3ZxX+vqgpO5UC43dDQYmsvGxxKOi+WkSlLkpepqooal5Q8aydsF7iEjOfOhYNDXtyrsoLruhulZf45bkjiOagtuwG8bTnQ8zxy4igKZGnWyUX2ILBsUDMfSCURhIEVmD9mPhBCwJEU+EdhBAFh1zymECiprCwb/85jyw1Tn3zfh1IKYbiWfWI1j7quoYU+yxh5DO1MeFmVVidYKWXH9ynA65gfEDWtKApyNjuRqsmpwRqLxhgs5gsAsDqKeZYjjqhyt1wucX9/f/TndTooZPFqCJpsBoMBwiAk1fEdhtiHgMm9vFhZUveZZRyeg9EGnu8hCMjuT0jiG7iua6V7tNbIs4dCnM/dM76vg8EAutZI09S+kFISabmqqxfxhfj7URRhNBohTVPKNopuli2ewjl308zPKqsSUnWEW9i4dnC3OovulkVpA0KbXe34+9RlaK1RGuJgqpI2fbwBbPviaqM7UVouSsoOP6m9+M7AHvOOcuyGmalMnu8h1KFVrWDZlL0yhoI4uEyhSVaJDYqEJOk0A2M3WE+hrmq70b6+vrYZeu7u7SraTX02E9pkYE+9ueC+gS9fvmA+n2O1Wm3Y2XYJDyhLW18HSLanLGlt2E4C7YtOB4UA7G5ZSYWqIiu9JElQlIXV6Wnvdg4Z9C/JUO2rDfWacBwHruOiP+iTxmKj9yalxOXlJeI4hhAC0+nUSn7sA07jJwmVL5IksS+oDQqrl3lE8kQUhiGCIMBkMkEv7lFG6Z0Fha+Bp+7fti4ii1kb1wAdiAkZWmvbPMLBIGtZfuI0sNmdRrSfNwZKKXiuZwPEXXOZkOLNgnIBYe0If6bnb5tAXBe+5yMIaTPuKGrGk1KSwkJJ78E+yxC/51VZIUkS5HmONEuJ5wZhg0Wtyff3JcerygoXFxcYjUa4u7ujtVK/L01ZrkScIiDkY7BLEEAVMs9d87Q5edK1oPA5XFxeIAxC+5yPxdFB4b4ncRDvpRHuvL+/h+9Raryu6ocP8AAds+0SnRXJ3bquc/N12uAXxXUpY1CUBaq8ZcwugF6vZ9Xw9z02l6Fu726pEafV+eq5HjXjJMmLJyjWgkqT1GYdz23E/h7B2cKqrqCc3fyy037gJlWhPZS2JXPyPEeRF5/P9JVhtEFlKqCiYI+5UJ72rGTRORd+5j2x89GxZdWugO+roxy4ngsY8p2HgeX5+r5PFIodAtFPgTXzirLAdDqFcpSVZ9KGZMZc10VVVihKaop4KiPsOA7yIsfV1RWKvEBRFAjDcIPi1JW17DHYczXrrOGpmkw4KwtBFoJaU6MGDOmmFmXRSb1CBlN0pKBNyuXlJZIkwXw2P8n8uzMoNMbQoGbbUk7pbut9HfCAnuPebafcmZMGwApYAvQibpdLtgONl2QO2zp/POh457C9697gzp05cyia/4qywHg8RpIk9nthGFpBTqXUfkLcTbq+LSLMOzbf962i+mK52ClnsA0pJPr9PuJejLu7O/uyMZn+PXGOTtX1dszPsTyN4zz00T05msvd3hBxhywLTtsO0xdkIs7J6zsJ1eTc2NJnq3VNunUFNYG5rrsOTkSL8/lGEkpFUWxs2I+9510KDJmXp5TCYrF4YO/JmUMpJUrzcsK/MAJG0MOpqsou+AY0f/f7fShHYTqd0sZLP03HcBwHg+EAw+EQk+kERV7AUY71D7cZsS6ncnm8ivX6cyxswgfUwNqLe9ZDOAxCChLzHPM5CYR3tZIlpIAuNbzQw7dfvgEA5vM5IPDzS9K8JdqlF6NfZkDfFWyXFYx/xO58R7BrQN1ZvufDUU03cpa9aDc1GA5wfX2NLMuwmC+gnDVB/hOHgbNzb9GJzF3jXLqsqgpFQdkHy29qJ+u335luvzo/BYxp7BDz2pbv2RaUpWxsEPDKr11Zrt1LfqZ3/FBq0kvQfi7tDRjTbsIwRFmUSNPUOno8ea5S4MuXL8jzHJPJhJ6J1tSJ7HtPuwZ1BO0yr4GBMuokSQQOhDn7anmWTfZwMBhAKTJrWK1WR1/Ha4C7yqMogu/7+HHzA4vlYr2hOHJN+CmCwlMEb1JIhHFoeVu1XmupdT041JoyN20pEIsTnbLruPAD6mZj3ovW+tkBWJUV0iTFfD6nhpiO3sNz4ZCFk4Mz13XfpFzInME8z21pkDO9wNML5ufzfhvws6iqhl4gldU59D0fjuu8SWDY7sTt+rx5aoh1av0kkIpK0k4j8J9n+YuyV2maoixL3M3uUBSFnSe4U7rLCcI2jKFmSs/17DUdezwhqLzvKAe+7yNNU1t2DcMQw9GQsr2NDFDXNjYc1BpjsFws7ZjgeKUTnMLXBnc3bnTPNi+fNNLyKwRITX+bY8hp+fbvrb9tt2cAgMuLS0gl8ePHD6DGWuZhqyS98btnRF7kcDJnY4HmUhGrnwP761Bt3yeWoQmDEHVdEwm6ftmObbVa2QBydDFCHMe2SaWLEjRtbN8zzrqcu0ON5WlY8PvYYLt9TRtyR83nVFVlRV554mmTsh/NoHyMWKBTMCDqT6UrKwdktIGrXatltr2Ra/O3ADz63DijYn9Hb46Vuq4fZAl/moCw6YBtS9C054C2AsSx85oABS5hQGVNmyVsnuX2eriNqqrw119/IcsyBEGA0XAEx3WwXC6R5dm6s/f8S9gGLIdQrP2PwyBEv9+3c9E253+fuZi1IKWU1t5uuVxiOp3an4miyMqvdRX8Hta6Rp3V9r6dKibpdFColCIPyB0vAS9InMFgte+NF3KLR7PrRRJC2OP3ej3EvRjf//q++TOtWfLcg4XPpda19YO0wV8zmfieT96yWXbQBLUtX+MHPgZ9srWbzqZI09Q6mTwHJu76vo+6rhFFEb7ffMd8Pu+8TMn2RoQ5Q6wdd86NAWfvANiGo0P4elJKS2jnBY0X/KoiCRzmIsFgo1PPbkR2PMftc+lCcHDoObQDnHO//8+B5zOG1hpZnqEoC3iuR5zDwKdMiGwtrLrF9X7BbRJCEOe8aUYqq9Ju/s69aXoNGFDQy/Iu2931rAm4Wq6O5qIJKeB5HuI4RhRHSNMUWZ6RxNMLGh452JGSxM+Vo7BcLjGbz6xUTheSGjsh1v9LUNd13Iut6DY7drTfxX3ea6UUoihCHMfWpIKbeRzXsTEFSxB1bRwLkEC8kNTAqWtKihlNTYj2546YbzsfFA6GAwAPF2ie/LI0w315j6zI9g4yjDYQSljSPpP4Pd8jI3e5zkIyn6ELO2CjDSpNqvbMLaOToiaTfr+PLMseEKEPgZQScRTbl2g+n9vjvkTvkF8urTWWyyX+8z//k7gapukA6yCX13JMxPq+clDInEjbWIHzELY5M9N+xg72Dwx5XLPgdF3XlGEqK8tRaWeQhBEvChp+VnRxoXgOLGfEwWFZlXbOU1LZppTndNr4OABVcByHbLW4+5wzOe/t/rwUnK3iQLh9nb7v2/mY7ccOhRBkqBDFZGu3XC5twL0PXURrjTzP8f37d0v56HKDifX3blUt+H++diWVDdCBl6/D7exoHMfwPR+T6cQG+VJIW5XsehXLGAPXcfHlyxfoWuN+cm97Ck7R3NXpoFBrjdVy9WimMAgCOC6JuCpFRNR9xrtylPWa9D3fynz0+30UOZXK2KKrqiprSn1OtAVheVJioVIhhO08nk6nJ+lE8jwPw+EQdV1be519dsJGGyuxsFwubYD46p2zx6AZb0opGxACsLpwACArCQ1tA6X3GhhyRrmua1RlZYPdbQcBDhx24onO1m3lgp8hYDhUdeGc4M+vqxpplZLElKPgOtSxrBxlF8XHwIsyQPMQd6B/hIDQwmAndysMyK+4KIujF2bXdRFFEWCIfpMmqXUiOQRZlqEqK7t2dMUmcxvcde37PjyfpM+CMICSCr1+D0IK2+RYluVe6xDznqUibcK6rm2zpDHGOm0B66Dw3Gv9Y/B94ghfjC5gYDCdTR/8zFPJCo6THvt+h1dmevkWi8VGxxG/kEzAdZRj+R77LsxxFOPy6hL9HnEWPM+DVBJfvnyhsmde4P7+nnYTO8bHtp3bW0MIsbEYO46Dfr+PWtdI0sR2jB46mTCvY5WsUBQF0jQFBGz270XnJza765jTISBezEt8a2xzhZQkWR8lle2Kc1xaQLc71Z/DqTNNxpAFEpu6a0dbIePHJn9uVNFaw2hjSyhcigB2d6E/di0CYoO7+9h5tv88BF2dpF+CLmUYuVtZF5QZ5swhi2A/5ZbDWZqqrKxIeZvT/BFgu2BNU0mJY7iei+VyiaIo1gmKPcGBizHke6xXlOkrq3VAuO87wO+nkN2dbxlshzoYDjAcDG2HsOM6cFxqmDKGgqDxeLx3mV4KyoTP53MIIZCsEltpcx0XgR8QFaIJOLs6plmqSCppvY5Zs7SsSrtx47V/15ixPMQd19jpoFAbvTYbxzqtzAuelGQrxOWuQwKzXtyD71MqeZWsrIaR67no9XpYLBdrn9EW7+bBonlCoudz2C4hGGPgui4uLi7Q6/WwWpELySk6ksqitErp9r89jieEsPetvdh0tYRh0WQEHNeBVNKKRnO5Wwpydqmr5h7vUUY+lA/z+Kmu3S5YNJidZ3Y1FWitNyY+pkUI+UgX8XNjW2D3750YpyiNHILtd+0UxzkbtrK6vHDw2OGy8s6FpMlMsxezNg/VBzpxja8Ifg/4ugM/wMXlhaXH1HUNz/P2Dljac2tZlJhMJuvsuj5OuJl5eF3NELZhQGsZS+dk+Vo+R0nqMSirEuPx+KDjV2WFyXQCKeRaqsd3LCd0uaLAnu95F2G0IXtbqVCiRK9H2sHsN17VlT3/p6gg7zJTCFCJl22E6rqG65C3L+9oq6pad8Xt+QxZ1DnLM/y4+UHHEuQzGUYhfvn2C4CW5EZH5ztda7iRi+FgiKqqMJ/PURblRpbwmJKXqdcE9EOaQ5iX2aVsyUvB56trbcdLu4uNS81duK52OVlArL1xd5zfXhnOraDvZ1/4n8KxzSpdhO0cbuS4cuRP/iywKY0BfLwxobVGGIa4uLygBpPVCmVRQil1UEau3UEqzFpX8iM7P62WKyyWC/vvOI4RhuHRiQ6jDSpQEkk5Cn7gIwgClFVJa2dZdvq+SykR+AEAwPVc/Pbrb4CgNSrLMvz9738n16MGj2YLH7m+TgeFSiqEYYirqyuy7slza7XG8gdVVdlFa9/sk9aaskBVhfliTuXBRs9JqtauqpVm7aQ9UBMQM99iuVzSbuEEg9paKhlsZGxf8lK2nwdnN2vTwc6Sl6DFa7WSLM1/h1AXXhN8nk+WD86UdftEd8HZg+fmjX2aHX5aGFqEtdZI0xTLBWUJbaLikE04WjI/zSP4qEE3QEmbtjYhy2KxEsJRaH5fKWU5ekyROrZR6ORorb0AlYpZUsd1XCilkBe57Y+4G99hMplY7uC+zYedDgoBIkbPZ3Ob7WCbIddx4Xou8ai0tlmsfR6mrtfcKtZ6q+saQgur/2ZbvtEd7+MHaALCu7s76i4sD+egbB52vUgwN8V+7wVBxUb6WtDgjMPYTqS+79vur67BgMqpruPa0lob3LWJen2dXZlIdurQ7Ti/jUaSA89939/ryj16a7yn6/58ps+DHbDm8zl1+WY0j7U7aI/JKu96Nw+pVgkIBGGAwA8wmU7s8bsIbmTiZsRdGVdO1tj1+NCh1ySSfN9Hr9eDlJKSKeVhAf1rop1w0Foj9mOEQYgkSXB/fw/XdVEUBX797VdAUKOSFBI16kebb5/ieHc2KOQgMC9yFOVaAoU7iPq9vu1G2sXfeMmDLUrSONwgzDcvM+vqcXfSdrTeFTCJuKqqjVT7xs8cuuA3L92GaO2hW7Qm0/bP//zPSFYJfv+v3zttOs4wMGvRWLTKZljrWHV1kgWefvm7Nvl94v3hI44hXiequkKVVJucW94Dn3CT1a5MHHK866trBGFAQc+Z9VWfglIKrueirmskSfJgffA8D1LIDVOGg2EazcIwQhiEqGpy3tJa2+pPl8DxieM4iHsxpJKYzWa4v7+HH/gAKFFRFqWNaR6VHzJ4tMkE6HBQaIwBBCyJn7+mjSZNqCarx8LVhwwQ13Fxe3tr07BVRfZQvu/D8zykWUoSAwce/y1gYGxWs6oqlEV5spfelkhlKyhsEVif/Ryz3jHz/2EYQtcavufb59tVsM6X1aza4q2eS6PwEHR1/O6Ln+U6PvF+YWCs+DdntU7RmLAR+MnWWN9awNtqDvx7Tx2Tu6Ndz4WBgS67FfAwWCamrsm/lytefH1xHAMA0iylXzigj4AhpUQURRgMSAc5WSXI8qyTPE7up5CKOt0HgwG01kiSxCaEAj+A4zjI8uxB9W3frHVng0KgCUC2pC6YUxiERLRsdx1va6I9B6uD2PodpRR8z4fnelglqw1rnS4NlDYcx8HFxQUEBG5vb5Fmqb2eY9TrudObNQU5EOfd5r4lav59tova7urs2oLfdg2xchHvJAj8xCc+8boYDoZwPRfTyRR5sbkQ77teMD8ZaOw0W7qgWmtAP8753GVLaisbjbxNJCIIQZmmNk+vC+tauzxuDDmKCCGs/zCDDSaO0WxkuK6Ly4tL+L6PVUINLewLfe77sQ2mKnBSpRf3kGYpsiyjNbWqoSJl748V9m43d+6xtO4VFLazPm8CscmvYM5BEAS244vthg55kG3Vcs5CCkMcDKUUkiTptIglQwiBOIoBAQQLCpaLsvGpVeLBLvYQzpDjOOj1eqjqCuPx2Aoc72xisDUUcj748uWL1e7SWsNzPfz6668kfFusFfsPObe3BF+X7/lwXfcoLaujuJ77LDYsa/FE0N3le35KvLfr3PWcD9W/e+rfn9gfUkn0+31rbVdVJNHDlZUN28AXoC111lZrGAwGUEphNp1RVWzH898udbrSxehyBN/zUZQF4jiGAJWRy6rEcrG0XsrtABJ4WqrktbBxTa1SfN3of3muh4vLCwRBgMViYTvljzlNx3XgBz5WqxXmi/mm+1e3YkKbmHIcB57noShIPznNUkrYCCDuxVBKIU3TzUqe2P9973Sm0L4grQyg4zoIggAwsDpDx0qvMHSt0e/30ev1oA21dz/FyeoKWFusKAqbiZNC2hKEFPKorl9+BqzZ5yjnxVy6wWCAL1++IPADlGWJIAhQVRU8z6NdYVngzz//RF3VneNxbINlaFzXhQBlPbvu3/yJ94vtLE6X56CPBhb6trZ2UsARjpX3MXq/7AywDsikWTeKua4Lz/OwdJZQlQLqh0HgLoxGIwoCy9IGfp7nQWuNXtzD7d0tBVjbrldHlGSPxXYWlBvmHNfBaDSCrrXl/W03Pu4L1t+tq9rGEQamc0oSQKOS0lhQcjA/m81sIOt7PqIoQlGSP7TRJE5/6HzR6aBwG65LWnxsEm6j4hNxAPzAx/X1NQI/wI/bH5av2HVwWzqr64dRSB3JBUnUFPXhHsjb/BXr5tHgOY9I3uHkRY7JZEK8hzSDkAK9Xg/XV9f466+/qPvbiM5yDDlb6vu+5bvUdb2hXdhldP38Xoqf5To+8b7hui5tjrVBv9dHWZVwXeKlz2fzDZ24Y6EkqW3ULgWfHMQwtt8J9qXOixy3P26hjbZqCa7rYjQcYbFcYLlcdpK2wxCCrEYH/QF838d0MsUqWcEYMkI4JltYlAXKadl5eSWb9TPktDKdTiGEQFVW1m0rCANEYYQkSWwi67nn+tR1v6ugMAgCXH+5RlEUmM/mGzcAOG7BEELgl2+/4GJ0geVqidvbW/u9ru/QpZLWDiiKIjiuA11rjO/HuPl+s/eL0y45bsA0wVErU1jhafNwIcheaTFfYDKZwHM9LJdLOC7ZahUFSehA0O47TdN9L//NoBR5ZbMEEF93lyeVT3ziE6cDawgqhzhcQRhgdDFClmVriS0DTKaTvdeNx/h9UpFPtarIZrOuavJdf+w4TfBX1zVm8xkWi4Wdu6IwstUaDhy6WqGp6xrD4RBfv31FkReYzqZWmP9YjrcQZEDAepNday5pg8cF8ym5C9n3ffKH9gOEUYjl7ZIadfQziRUBm8XetXZ1OygUlAVzHRfD4RCD4QB5luN+cm93DKd6kAYG88Ucvu/j5scN2YWJbtoCcQMIe0OyzY0xVCIAAEgqIdzf35NV0J63yfM9fLn+Yi3QAj+AVBJGG/z222+QUmKxXODu7g5Jkjx6HCHIWYODvTRLYUBkYuUoW47OTd7pgNAYQ+KpeWH/3eVd9ic+8YnToc2n5y5QIamyUeQFqrqCoxxEYQTlPO4d/dixYYAwDtHv9RFGobVdcxzagF9dXUFKiSRJcHNzgyp9OhOZ5zlJq2hNdpdCIs9z4ijKteuKVBK66k5Q2J5PBSgjNh6Pkee0PrBkDNDKojWL217rtYGVtum6QHh7s8CNn2xVKoTA5dUlVssVJvdra8TtJs590OmgkHcEcS/GL7/+gmSVYHw/xmJOXIiTasQZ2pnc/LjpdHACYGOycF3Xdkrf399Te3oQ4Nu3b/B9aojYt8OMA8G8yO3OGD49j6Iq7P1ZrVabBN1HzpV5Mdk4s5lDDgaLonh+Z9MFGGyQx7ddXj7xiU/83Ghr2AZBgLqqMZ1NsVwu4Xkerq+vEUYhXMfd88DrP7XWKHKqnnieB8/1UFWVVZTI8/xZfVejDTyXkgN1RU0ZQlGTpqMooKh1TYGheBg0dCE4EqBMXlEWuB/fW167FbY+skrD2dGuZgefQltZ5OLiAr7nYzqdYrVabSQqfkpOYV3XSNKEdlFBiMVyQR3HTVNCuwnk2NKxMSRSnGXZOtvWYfBOr9frIe7FmE6nyDMS+jaG7JKKvNhb6JPvg1IK0+kUnutRc4XnIpABlYIXC9s5/BwHsCxLTO4n9mdZZoBlhdIkpVJsTc0xXS1ltGFLDeefOz/xgdCFxfrUeC/XpKRCrWn+iqMYjnKQZimSVYI8y0ka7ZLWo71dmprmjqqqkKZrqZEwCoGI5tDFYrFuqtRPS6RVdYXlamn/zhklx3GgHEWi21WFqq4euB91BQZUDRMQVkmDmy22VUP2HUOPlZzbEi5dazZpg7uvL64u8Osvv8JxHCwWCyRpAketQ7rnOIWPZVY7HRRKKREGIbI8w59//Ulk2x0B4Sk/T+umc7fDWSB22Ih7MaIwwmq5wu2PWxtAB0Mq9U6n00dlDJ6CNhp1VSNNU4RhCMdx6DN9Y1XSy2otLPrU8ZeLJZJVYkvbVVlBKgnP8xAEAWbTmdXNUlJ1Tg5gG13mnnziE594HbR9iYMwgAF1guZFjlrX8HyPdOKq+iA+IQR5/RYlafSxVZnjUDOL0dRowHasT6Guavz1559AU5UpyxKu49rSo9Hr5sEuz2VsmsBSdNroZxsb9/6M9voluqHb+Bzqukav18PV1RU838NivsAqWdGGQR5/7p0OCjlrJAR1XPGOp41j08fclRV4Af71X/8Vt7e3uJ/cA2L9M13jFiqp4IUerq6u0Ov3MJ1OyQqQx7akl8hos9s/8onrsXI2ghTkHUVk6jAMaXes07V4KH/ejmdgicANQZZFNgGaiIIggDEGs9nMnlOXX0bP9xDHMbIsQ5qm9tq6vKP8xPvHMdygXcc4BK/xXm5zx3iz2dU5wBjyQo/iCHEcY7FYYLFY2E03N50kSYIwCLFKVi8+thVpNhTQSSnh96hEzeoXLCtT1uWjpdP2vF4UpQ1wWLB6dDFCGIaY3E+IZ95xCCHw22+/Ea3r+81aXoc1hQ8c1wLU1awUZU25YSMv8g2eYRey2PwM2+fiui6ur68x6A+QpRn++v4XsiyjjuwdlbZH1+dHOpA7HRS+FZg8rBQFiFJKCqqawWdFSTswSIB1sBrHMaqywmJOpQUOBlkTMMv2f/GFaGztGkgp4ToudK1RS+Kh6FrvLc7KcFwHeZ5jdDGy59i1oHsXuPziKIcymoAtZXwGhp/4xM8Nngd9j3xmda3tYi2lpK8boKzKoykwShH3r67rtXZew5/fV0dPCIHAD1DrGlEYwXEcLFfLjQ16V8EBreu61NSja3u/hTmua7quKSvr+z76vT7xF5vO5nNqNb4EcRxjOBhCCIHJdIL5fH7S5/hug0J+eIfejDZ/jWVWlKNsYwQTWkW93pmwYOa5g0OlFOq6xt3dHXzfR5qltMNspAvCKERZlUjSxHIzDh3kSpEXNE92ta6PEsYUQuD6+hrD4RB//PcfyPJ1UNhlPiGLVldVBcddi9RKyJMGhnwvupw1+cR5cO5559TgZoLmH5R958xYI5XSlXfAGGPLu9PpFEmSWI6067rWl3fDK/1AsE9xWZVQhsrFRpuD74cxBhcXF7i4uMBquaJzbwKsrtzfXXBd15bkfc+nxESjDXuMcHUbjmrMMIAN948uv2ur1Qp//vknjDGWa3pKvKugsJ3uPIUPLZcEhBDoD/qQQsJzPXieZzOFlqir1+XCc2cOq6oCDGzplZs9WK9QCEFdvVV9sJ4TX5/jOFBKEdel9SIeeu/jKMavv/yKNElxf3/f+SzhhhSFoGyB67ow2kAKiaome6tDbke7LNCFzcYnPvGmEOs/rcpBB18BATq3Ii8wKSckpSWl7d51XNKM04a80g9ZpHk+VVJZCZmiKuzcw5vEQ+RTDAy+XH+B4zqY/DnpbJawPdcaYxCGIaSUSMsUQRhYi7csz2hNrvdb19rzrVLK8kCtvBjExud3FVVVEcUNjcvWiRs0Ox0U8sXaBymVFeVkNfNjFlK2j9FakwWQ0bi+vsbV9ZU9/vh+jL/++gtGEIeuC4s37645GGwP6tFwBM/1Nngje5UbmgmQvY57vR5WCXlMcyMI37OnXhxr2cSZr+Znr66uEIQBfv/H7xu/37UsIQfA2mi4DknqGBirH1bXtfWanC/mezmxtHejG6bvAmsHnWaB7PLk9IlPHArOEm68C4oaIaqyIh6yOX7jfwpYHTy1nneZe+a6LnzfRxRHmM1mmM/nD63jXnB8FiTu9/uIoghZnlF5M/DtnLuLX9bGNgeef/brl68Iw3CDA9lFtINCJRXCgJocLy4uMBqNiHcOg+l0iv/+7/+m9RsvSyoYQ5aqgR8AgtzLlFTWCYwbiJgCkGUZjcEO7FKeijdOnSUEOh4UbqPWNXSubanhFOAdied5KMsSSZnQC+o6EBDwPQoC8jzfaPfuErj83e/30ev3UJQF0iw9KHAWQsDzPLge6R+WZYnlcknZMX8tE3Ao8iLHzfcbTGdTG0h1LSAEWguBlHZHWVUV6orKFywe3vzwi8ABIHM222Rfnqg19LuwVvzEJw6FFNJWaIAd89P51+FnwRu6OIpxdXUFow2SVYKyOJBTaNZUHaONNQSoqmrv+dY2Czao6xp34ztMJ1PMZjMb3HYN7YqM75Ofr6Mcks5pqjJs1hCFERbV4sUBrhACQRDA931cXV7ZxEq7usZe0atkZTcmHxHdjHIegeM41qKnqqqdnbX7gHmDcRTDdV3cfL/BfDGHlBKj0QiXF5cbzhXtl/2cGcN2FotfJNd1MRgM4LouZrMZ8mzNbVFiP4V9rTVpNuYZqrJCURQIggBSyv13wVs72x8/fsBxnGdFr7sC5pywhdUqWcFoyhiyQOxLwYHmUxkQIYRdFLu6o//EJw6F3RhtBYQPxnrHA0MlldUSHPQHyIscSZpYSZm9NuINP74sS6xWK1pram2TFc+JVe8C+x0DZLnHHcie71kJsK7BjgUYBGGAIAiQpim+33xHnueIoxi//fYbuWsdoK9oNDUGFmVhFTYiNwIAlEVpu4/LsrQUsY+ITgeFzKPg9G4Yhri+vsZivsB8MbdBIZcqDwnUHEV+wTDYlL1pdm55QcEVNxl0CdyJJaVEFEeIoghFQY4jta4pSyj332UabYCSNAa10RQANZ6/rE/40uxYrWtryyOlRLJKyA2gXneSdRF8jcojyoKUElVFATKXjtt8n5fwoSwnaEvuiLOHLx27Xee8vBbOTdv4xOHYCAJbhH6bFX9nVAnO6g36A1R1ZUuzB6EZ1uwDzxqunu/ZdWefMuEGV1lS4iNLMxgYKKks/WfnqZz5HWNaQRAEEEJgsVwgWSUUzLkFirJYV8L2CNy4fGxgcHNzA9dx4bikJBGEAbI8w3g87mzA3AZbF2q9Tgrx31nk+xh0OiiEodZ/JcnMOwxCBH6AlSINKOUoUpJvWY9ZXsILBotSCtfX1+j1e5jNZlitVnCd5iU0mgIgvZYdaAeFXekOZU7LxegCfuDbzriqqg4qswsI63Fcm3WHWlEUKFEiz0ms9aVcH11rwFnLC8RxjDRNN3iJ556IHgNzCD2XRLeLvLDemyxfxHhpdqBNFrc6h4c8p47es0/8fDj1WNvWXrRzwDsa0o7r2I7e+WKO8XhsnUj2vV/MB+fsI0Al3+ViibIoKRDKixfNldtrEicNSpQbPPAuzh9CCChHIQojDAYDGGOwXCxR69pa9DmOgzzL19SdPY7tuq69/qquEIah1Sjk43GX9/b9eWlM8RZoxzi+70MIgTRN4bkelsVy57nvg04HhUIIuJ5rB4Ql22pjuRYb3bVNtualDy+KaPABwHK5JFNzkDSN4zjQtbZlzk5lCbd0lC4uLjAYDpBlGZbLpZVFOGSC2lXWybIMeZavg+89gmF+XkIIxFGML1++4G58h/lsToLbHYWUEmEYotfvkbZikaOqK5tBZs6p5Z288Da376vNEnZksvnEJ14T7e7O957tvri4wOXVJdI0tRvxYza4Bo0SRiPLUxYlSlHaysQ+/vDtIFtKiX/553/BdDYlk4OO03aUUugP+giCgNbkqrKScMz92zdzugvc2KQU2Re+hwwhg8eYlMRplUpSAxHINezYe9PpoFBKiV6fOmAd5ZBBuO+h3+/blGmSJCjLkhbnPd9HzvaslitM7ieoqgoykHClaxsL8oK6tU7ppnIStAJD13FRFiXu7u6wWCxQFC/bVe7zOVzGh8CzncdtSCVtF3K/30fci3E/WRucdxXt0nyRF1itVjRBwUA5Cq7jwqDZnPDGZM9FzjadHNlF/4lPdB3b1J52xtz+uwOdxi+FlLQQ393dYTFfWDrMMbD3wKwTGxUOS0a0O3l7/R7yPMdCLSyNp4vQWpMNanNv7+/vUVYlrT/awPM9kuo5UPanLc3G5f+8yA9KnpwT7FYmFcVHF6MLS1+oquP9rLsfFMY9fLn+YgcB8+dYw2h8P8bkfrJXoMKoKxKATlOyboMgjlfgB3BdF0VBaftjG1peC7yrnM1nmE6ps8wKcuP4DBT7fXIX8yFlTmMaHouS8AMfZUElebYZMsYgz/O173RHJizeCCzmC5RVuSHlwOUGrUlM1ZaDW4vac/eJyeXtbuRPfOKnhcC6mtOaTtuuII5y1nxlc7gW6ltgOp1iuVxiPp/bjeEpsGsuYezDOQawllprGgdhQM4rAhuJjlPoz54Ehsq6TOWaz+d2Xfc8D2EY0npR5AetyWwVCNB98FwPWZpRsNkYPLSrYV0KFNtmHVJK+55woowdd5RSNrt6KDodFDLfCgDG4/FGNtBRDobDIfEE+Of2vA9pmiJNUzqe45BNnFLo9XvwXA+z2QxFWZCyfBMEdALc1CCIe3I/vn/w/VMMaJ4sOFBr6yG+FFprCFfYZo26rhH3YoRh2JwqEX+11tTZ3I2Y0AarTB7nydM63kiBPMspKNxh+ffc/efjsbRNW3PyE5/42WDH9VZDiRXJd8nOjDs/u/4eLBYL+/dTBg+7urH3lRTjjFhd1xgOh1CSsmKji5Gdg8uixPh+vPP4Z7v3zdhgUwa2EXUUaeaGYYgkSZAm6brStMepSiGtBE3ci6E19Q14vmdtCzc4rh2AQKsJ0QBGGOuoxQkbKUnCByCBdSXJ0/lQdDooBEBK8kWB2WyG5YpIlEop2511SiilAAFLSE1Wif1eZwLCLbz6C7wj2N5nN8k8kCAIbEDluq79vlIKuta4G9+hlt3VheKuYddxrZZYkVM3W9sucR9YftUnp/ATHwS75iue07mx0Gizl8JBV9CZjJsgGTLu4jUwGI1GGGIIgNayxXyBxXKBsugOl257/uQNs+/7iGMK4lbLlaV07QsDA9d1MRwNEQYh5os5qrKySZROlpFF0/wCbe0UwzCkREJFftZSSgwGA+L99w3u7u6e7DB/Dt0PChsYY8i2rcnmOY5jeX8HHY+5G61BoLVGFEVwXRfL5ZK6yUBimuwV2ZVB82AC6igvzXVcaKMR+AGUVMiybKMDbtAfIAxDCFBTUacaelrg3aPjOJCKOtGtPM8JsE2873qm5BOfOAkEbCZEG22zhPzfe8EuzuS5YIyBUAKeT4odWZYhz3MIkGtH4Ae2mdK6g9lfPttpPwAHhUEQoNfrUQ9Bmhy8RrSfUV7kyLJsrYAhKSMnhYRGdxJAxlDGt65r+L6Py4tLDAYD+L6PoigQRRGqusLV5ZVtyJnP58izA+WR0PGgkOvoNiCTwrqK8IBhEetdreRPZWA4TSyxFlP1fR+j4Qhaa0ymE/u5XU7k8EAASBT51IHr0Vmshofo+z7xRaYzlFWJqqow6A8QxzF1IQvAVd0NCnl8hFEIIQSKsng4oe4BljTi8rNy1Lp8IVo8zk984ieGFNJmCdv83K6Dz5NFkLuU7edSI5sy3N3dYb6YAwboD/q4vrreUKfo4j1nnqnv+ej3+/A9H9PZlPQWmcJ0wGnXdY3FgpxQqopkaYQQqMomjujQpMtjylHkha1rCvjKsrTSPZ7nAQJYJSurs8y8yUPjgE4HhVpr2/VZ1zVNIM3iaZsUstxmbHap4j/2snL3cm1qeK4HxyWOou/7JJiZJPZn2p1cXYTAepcN0CB6DZ7LIeAXj5tMsjyjBp6iwMXownaTdR2O46Df66Pf7yPPchRFsUHoPUSbjIXCOQPJx+GAsUsT1Cc+cWpwQMge95af+w5KxxxMtQWUuzLnSiHheR56vd6GsLaU685dXlOZt9cpZQ2skz5RHGE4HKIsS0ynU+J4H9iExNVG1jZ2HOKx1nWNLMus5Fhn0IpfuKdhMplgNptBCIF/+ts/IYqpfHw/vkeaptaJ7JhNSqeDwrquMZ1OoaSiBRQ0gH3fRxzF9DDzzAoK7wNOJetaQ0iBfr+Pfq9PHaeLtaciE1DP/ZI8Bt5RmcrYppsueedKSVI0ruNitVpZ+SApJRy35Sfc4SwBcyI5S5hlGZUemp3lUdpkDaewLTbeVf7qJz4euFoDnLYkykLFyiFZsLqq1w5VHS8db5D/Adu80T7lXQ0jb4nBYIAoimyzJLtgsJRWnudWm29bm/bcEEJYe9FBfwDP9fDj9gdWq9VR93O7wYk1eLm8vqthsKtgaoAQpJVbViXKqrQ2tMdcR6eDQoCyhbrWkIo044w28FyPLN3KVrZG7D+olVKUipUK/V4ffuDj/v4eq9Vq/dmHmJu/MaSkDCpzDbZFSq0URIO3fPkH/QEG/QG00ZhOpihyKhUrpcgppOHmnUJf6bXAWULP9bBYEEGby9xH38umo6yq18b3XQ2OP/Ex8RoNFLzws7xGret11/E7GP5CCHiehyiM4Ac+xnfjTSkQs876vzUcx0G/34dUEqvVygasLLoPkNdvVVXwXG9z3j2zFBBz+IMgwPXVNaIosvI0p6QWaaNRl/W6Ylh3uMmxtX7zeuN5HvzAt0FhXdH/x3QdMzodFNrOTLHmbgDkROJ5tEAfM1CUUrYmb4yhBb8RIuV2767sntpoW+y1d3m9fg9BECDLMst5Y+2vjRd9u8r+itfo+z4MDJFfi9zKCsVRDKUUsjwjGQp9WAfvW8GAdL3YMQY4zbnaF35rMn4vjkSL6wAAMRlJREFUO9ZP/LzY7oy3shg75p+9j93M61pru/GH6e6GiPnDLGgvDGU3/cDHxcWF9Ymvq3qdSDjTpXieh1pTlW2xWFh+cl1Rs4KuqXwsBRkLbAT94rxBOc977OCSZRnu7u6s3V1bhuaY+ZcpV13lsAM7NCubd68ua/R7fdu4yRurU1EBOh0UbkMIgcCnTqQ8z0ncsj4ucFOK/JMXiwXKskSapnai6uoEBVCQLCSVjlmo2vd9m1K2fppKQVdb17J1u16TJL1YLlCUhe30AiizGYQBACBZJdRV3pRN9/W0fAtorbFcLpGIBEVe0AZF4qTlhs8g8BNdwrb4fbsh4RTzIjdZwbQCw45WZdiXmIMoXnxr1HAcB2EYwvM9m+2varJhO8c7LYRAWZUY341RFIX1Y5aKqkmOcpAk1MErleykMYM2GlmWYTwmHcXlcmnHxnYJ+GAIrEWgO4wNa1lBbiZ+6GMwHFD8YzT6vf76509AdXtXQaHruhiNRvA8D3djsnTjHcUhRH/eJdRVjdl8RrspTdyWXabYXQGTcNs7A8dx7L+tM4jAhk/kOa4nSRIiwJZUWnEc4ooEAQWFy9VyLUrevfkJAGUJVqsVTa5CWg2oz0DuEx8BrMDAPKxTzCOcVbM6bB0NCIEWx1EAEtIuztaJyOpyr+/TucD8ZC6Her6HPM/hKhfDAekULlfrrFttqIHzKSeVtwavzfPF3I4NTn50eZy8FtqBaxzFuLq6glIKd+M7DIfDk6/r7yoo9H0fw+EQi+WCrO2OGCDtbmWtte3OgkGnA0KGUgphECIIA9JsVA56cQ9CCFxdX2E4GiLPckxnU+j8jC8Sj+dGBFsIAd/zSVTVkPF728C9q009nMVkOZquZjU/8YnXQNs39lTgDe17WOilJCeMKCKLVd/zobXGaDiCHwQYDKghoqorVFWFyWRyliyUNhq6ovuqpEKlK5sk6PVpfeAOZO707pIuH4MtXLVZ0wvazT0fEVJKjEYjXFxcUAUuL+A6ayOIU9mlvqugsKoq3E+oEYQX5oPRBCnGkLE0gKN5Mm8FYwykoJf8+ura2qS5rgvlKLgeDZTlggS4q7KyGVXgba9vo7NNAlJJ9Ad9+L6Pu7s7ZHm2/tkOv/RcPuMddlebYj7xiVPjgeVai/96LK/ryWOcuemhDU4i9Ht9XFxe2IoB3Q+DX3/51ZZl7yf3mEwmZzlPXhOVokymEgpFTiLHnutZBQittV0TurgRt7zVdlLhud/ZIwjfd1yds8zc7nIvygKL5QI3Nze2/F1VlU1khUGIvDhcuBp4Z0FhnufkN6sPFw1uo2svwj5olzRhgDAMMRqNUNc1JpMJ8jxHVVJn7zbesrzRbnJhmx7P81DkBXFFOt5g0kY7u/wezvcTn3gLHDufPPb75256aIM5z6vVisqZjRbgcDRErWuM78aYzWcwxmC5WJ4tiLCb8EZyTSmFOI4tD5/pOuemFb0Eu5opn/z5Vx4s596g6JrG33Q6RVmU+PbtGzzfoyRREyAWRXG02ca7Cgq3G0C2yc/HDu728br6ojCqqsJ8PsdysYRSCt++fQNAUgPj8RiLxcJOZJxZPAe45R8AaUH2+5BSYrFcIMuyZ377E5/4xDlgM4F4mL3f7ko+BufW83sxGq7gfDHHcrWE67joD/oYXYxgNClXjMdjsl4tu9PRKoTAxeUF4ijGYrHAfDa32rv8feD9VMk+MrgBpyxLa/3nOA5tQrSxmUTP8476nM4HhW0ui+u6lGUqCuR5fnKR3+2gsKsTlTEGtakhtIAW2vJcgLUloNZ6o7kDWE/0bxkgMm9IKYXhYIgoipCkCXVOfYo0f+IT3YXBRtbh1ebDhsrTZTDNqKoqy3/u9/p2493+vygKKOd8fGMpySFGSTqHwWBACgqrJZI0eTLw62Ip+RNr1BXRxPI8x82PGziOg7Iokec5/MA/OiAE3kFQyN1pUkl8+/YNvu/jzz/+RCnLo4IKtlZqvwCOcvDlly+o6xp3d3cPdOO22+Hbv/uWtmQsNWNAsg5sbs5/ckmZ74/WeoOE+tbEbkeRmGrci1EUheU6sqL+e4Hneri+vgYEcHt7++7O/xOf2AuNbAewKeR/6kyh53kIggBJkth3iiW1eHN+bkFl9sflzt7BYIBev0fNZmItl1YUxdn5Z0oqlFUJqST+6Z/+CUYbzOYzJEli3cGAtSRLl4NAKSS+fvuKwA/w4/YH0jQF8HEzmtpomIpikfl8Tu9H05BTJ6cR4O58UMgaUa7jIggC262m65b0yqk+S2550HY0Uwisd65BEODi4gJCCCyXDV+kJOKpbaA5o6OJEM2EWlVYLpZYrVZIkqTT93YX2JbL8z07Jkt8BoWf+DnBzhK2+UsApt7hL3+Kz2r0Vs+o5PIk2I6SteI8z8OgP4AxBmmaQkjSJjRovJBP1AV6MFofXxYlkiTBdDalsvY7yMoyWF/R8zz4vm/X+lNuSt4j2pS5bRWVU6DzQSEbVwdBAEc5WCwXqKsajuuQZ+YJ7WlssCTWwYz93itIMhyDWlOGcDQaYTAYYLVcbRBOuXRw7hIt38M8z3F7e7s2vm/Osd0V3WVIKeE6LlyXOrvPPvF/4hOvCCEbwWOpqBwpmqrDKcWORfM5jVvVe8j+MA2m1+uRF682iON4Y4E+93XoWsNRDnStMZvNsEpWa57jlhvIuc/1KSil4Lo05zquQ5uUDx4QvgU6HxRy67/rrTOFruMi7sWoygrj8Rjz+RxZlnUqaHttSCHhez76vb7tRO73+1COWkslnBH25TWwxOayKB/wGvnPrmmV8fm3S2b23uJTkuYTPy/YzYQ3mY7roK5qKxHS3mhul3bP1dD26jB0ba7nIoojGBjMpjMEYYDr6Hoji3XW02x0B5WgMvFiuTipE81bQgoJRzn2f557PzLeYtPR+aCQeXOOcuB6LsIoxOXVpW2rhwCyPFsLcu4RGIZBiCiO4CgHZVVCKWVFleurGnVdWxJnWW1yGHd15b0VDCjLNhwN4Xke7sf3WCwW8HwPTu1YY/lzdpTxYiGF3JkNZFmHrgWDbQRBgOFwSG4xMBj0B4h7MdI0xWg0QhzHJBOQrFDk5+USfeITp4AxxpaMHYfmXCkkpCstiV0IYbNP29SU7fd5O0iUSpLYvkOLvKMc8uqta8stzLIMWZahruvObL7KqoTruLi6usLFxQUpP6xI+SFLSUWhC53UbT3VKqs2zqvrEELAcz1EcYQ4iqGUgud5iKIIrufi27dvuLy8RFWT8ob1df5g4PeC+aGnprp1PigUENYWbbVaYblcUrbQdW3HLbC2YtonWTgYDBDFEVzHRVmVCMOQSJuNUr1SCtPpFEmSIMsyWzo8N4wxcD0Xvu8jzVJ7TzzPg+u4tvsMOP+E8FTQ1+WAEIbKF9fX1+j1enaHVlUVenEP/X4fRVFgNpuhKAsUeXHuM/7EJ06Hppxb1zVqrDd1SqoNJ5/25hN4er7hRV8pReVAKWH0+ncdx0EYhHDdZm5LU+T5cUK8p4LneXBdl7yFixKL+QJSSIRRiDAKN6lGHQjC3uMGVQgB13NxeXGJr1+/wvd9FGVhuZBXV1dwXBfLxQLz+fxdXuOxUJICZb52JRR0rVHVp5NB6nxQCAFEUYRev4flYonb21vL41Bfjmv7n0xJ5JnLI0oqVFWFLKfOWM5GSkkNHW2NxHNjuVzi7//5d3ieB6kkLi4u4Hs+nXdT6mlzDD+xH4Sk0vGPHz/w4/YHYGD5m/P5HOPxmITBDT5kFzKX18/dGfqJ1wE/WzuXsG6hS8oHh5TxjDEoygJKk3KCoxwbYAohUOYlVsuVtTYz2pw8C3IoqqoiYWAA0+kURV7g6uoKcRTbRMJHzFqdEsYYlGWJu/EdlqslpJTwfR+D/gB+4OP3//odaZrCaINk9f6aFY8FvwvsYOb7Pq6vr/HnH3+i1vXOyuAh96jzQaEQAmEYIggCTO4nMJoGDptk84u4XcZ4CZJVQvZwjgttNEajEfyAAqvxfIy6qm0pls/l3GA5GjgADFAUBeJejDiOAQGsVisqq6Mb5/sYWHKiqxQRYwyKvMBfi7/gui76/b6V9ql1bcW3pZQoi/LDWN/Zd4Gf3TvqZvzE8xBCWEI/z69VVVkqCI4olhhjkCSJ1VZzXJKq0kZbmhAHXrwAcvB57o0Hq1LAAFVJiYIojgABLFdLUnzoUNLgMXShEWYXjKHAOk1TFEWBJCE9xW9fvyEIAhuUT6dTa+nalQ3DW0EIanbN8xxGGwyHQ/z666+YzWYop08nJrbv03bnchudDgqllBgOhhj0B8izHJPJhBZiJa0gMnMJAVDJw7y8SzgIA5vliaIIvV4PRVFQ2aSikgl3xnHQee4XysBYQWjm/qRpiv/4j/+w56ZrbbunuzYJ6FojiiMsl0vAAI7bzSHI0j7KUZZfNRgO1t3HzeJZ17UNjgzMQRmU9wQ7iYh1thBic9L5zB6+X/CmM4xC8lUtKxJtLivAgfVVN8ZsbJhfdOyG4mKMoXJX86rw4sQBof0adi9a5wCrXGitrVTP77//bt+BoihO4gd9CuxyoGlj+56e+3z5HOz6pTXyPCcHrEEfjusgTVNkabZhxvARwM9KCmkbneq6Rq3rpqFUIgojLOYLuK4LYwyyfO0Udkjg3Om7q5TCxcUFXNfFeDxGkibUZKEUfM+HEAJFXmx0xu0LKYj47Ps+kZubNOz2zexkVmvbMN7wH61sDs6/y24jjEJcXV3B9/2NrGbX4CgHaNgJUlAZQwppxWnZNYb//tGkEli7jS/ZXrvZ3IV2aex94uXgDGFVVVTGbTRcjTFWUmrfxaYtmqwk8Qo3ApJ38voYY2Bqs5alMuvFtytBbBuu6+L66hp1XWN8P+483UUpBSXJsxnAWhCcxdQNBekfbm5pkg9SSmtUkWUpal1b6Z7HOLi7MoWPcfo7HRQyx2CVrHA3vrMlB9YtFKAsmQ0s9ixlsV8gi2MmabJ2OpECpu72oONAuNlTb3yPF+mupdi5FFtXNWULOwqDNR8ziiOMRiPq6Gs4plJKm8mQ4uNIJbTLelJKK5DO4DKQ0evAsNMNRZ/YAAswM5+aSf5cmQFoQdZG770Jl0Kiqit4rgc/8G3W3W6s3sE71N7omGpdhenSHLsN13ERRRGqqiKljY4GhTwOXMeF55NAuIBAnuWWH8+SSB8lINy23vV9H9dX1/ADH77vw3EcXF9fYzAYwPM8zGYz/PHff9jfP2Tu7XRQWNUVbm5u4PkecVFcx7pJOI6DuvGZ5J3rvjDGQDkKgR9AKYXVagXf9wF0I6X+HDgoafO82iWMc0+021zM9m5aG42yLNedjNtZzzODMyK+72M0HMF1XKxWK5vl6GpW4C3QfjfaNmhtIjQUBQ9Mw/jE+4HW9G5WVWU3PVJKW7azQf8B7yvTXhzHgeu6Vl7jnBJfh8C+/1v+0F2A1o3vcXNe7Nlc1/XaoaaDsCVkQXJgTO8SmtZ8GFj+6UdFv9fHcDi0G7c8z6ms7LiIo/gkKhidDgq5kaIoChvcSCWtm8liMSfSZZO52LdcJaVEGITo9XtIkgR5npPMjVkP0C4v/BsBHzsCGKzLyB0o3/F9dB0XyiG7QuaFeJ5ns3HthaYr91wpheFwiKurK6xWK0zuJ/jy5cuDYLxL5/za2OVFWxYlirKwVAzmndmMUoOu8Vs/sRvcdSwgIB25zt54ng0uDs3+Mg2DNxNpmtomufcyNngctzUYuyIBBtB7FwQBXNdFWZRk/uCSVJlSCp7rWS/rLnVMO8oBREMbG5F163Q6RRzHiKKIfuhjTLNPoixLfP/+HUVZ2PFW5AX+7d/+baNyYzPaPxOncBtGG0hXYjQawfM8zGfzo1LhnudhNBrBGGO1/qSQ0OjOi/IcuEuQG2FskNWBkp0QAr1ez2p8KUmt9HVdI/ADXF9do6orFHlBMkB1efYg1qLRKRz0B9BG435yj+VyicFw8KGIzttoc2t3ZaJPJYvwluiaheU5wW4mFma9EQdgg8JDn6kxBr1BD0opJEmy/twWP/U9wPKJt96HLmA0GqHX65H+blnaTZqUEoPBAEVRIM9ypFlK2cOOnLc2GoEf4Nu3b+gP+hiPx1gul4iiCEoq2337CbK5TRKS5fF9H8pRUI5Clq2bTA6tZr2r1U1KiTiOMRgMUJYl+SA3XWGHZMWqmia4JCVpmve62Btj4PkkXJ3neac4I77v0661EdUWkrhJylWWPLySKxRlYdXZuwDu8s7yDPWktvQFJQ/TaPtp0HT4A5sLeVee2yHYtjT8yNhuUtNGwwHxuGFAMl1HSK/oWtvO/jRN4TouVWbe0TvFagTtMX9MoHxqhEFo51zHcRBGIaqygpACw+EQZVliPp8jL0jaRKiO3HuzzlJPp1NMp1NyMnNdyoB15DS7hLqqUTvkBuQox4pYH5olBN5JUMhSH0EY4PLyEgBoUGetTpsD9NLYkSIvcpJhaBxSmOdSmerBJNkFWHmchh+ia40ojDAYDHB7e0s8DObxnXmxWywWyNLMGpr3B327KMwX840ux319U19z18hl0vvxPWVjlcTl5SX8wEeWZp0qu5wLWmugbgUSzU6+3ZHdZbTldT5BYJ4cd9YqqeD5HjzPQ1mWKKvy8CwhDIymqozWmuatKILjOFb8eZeaQpfA45qbHeMoRpImWCwW68Cw4Rmea/xzwKekQlVX6Bd99OIeyrLE/f29TRxUVfWgUeycMCAJpPF4TNI/UuLq+gq9uNe5Uvdbg+fVqqqQpInlcEspUZYler0epCLNXODwLCHwDoJCniQc18GgP0Av7mG1WmE+n2946h4ivyKFtCUMXWuEYYgiL5CkyVpao3W8Li1ybbFuKcluaTAcYL6gCQFozl8/3DG85XXkeY6qrOBU5F5w6VwCAkiTFGmabjQi7H1er9icIiBgtLHp+DiO4SgHWZbR2Ks/aAMF325BpURRb2YNuWFgu2uua+BJ8ykNty6e91tAGw1hhM0yMYViMV+s5UEOAP8e6xE6jgPPJT/lNE2JJN/RW74tT1YWtBB/+/YNf/71J5aL5Vqz84zRrICwwTtAY3jQH9gMXJZlWK1WZzu/51DXNdI0BUDNJlJI5EWOZJV0qgL2lmjrN66SFZI0IcWVZvOmtbb6n1mWHT3+uh8UGgPXdTEcDHF5eYmyKnF3d4dklZyc/zeZTKwMQ1VXZ325XwJe2Nh5gCdsJZXdWWhoiPp8XAzmOAoh0It773ahzfMc32++23v+YYNCYOfCzVle5Sjradv1e9TOaHal9NcVGJC/ehiEqHWN1YooHqecRuq6xmKx2DAh6FLmqo22ckJtajjKQV3XVJUBdVRLSMtP1fWZumQbHbuqqkiKJo7g+V6ndRQttjq5y7LEjx8/gB+0UeEs2EcEJ3hYh5Az7QDgBz7CMESWZhQUtnRiD0Gng0J+qTzPw3A0RBzHuLm5sRPUA2P2I1/CNEmtOwN38nYxMORA0Pd8+IEPpRSiMILnedTJZ2BLsrUgDtC5LkMphbKkDrhebx0UtjUW2+hSmb6NoiwszUAp9aFLGe1ntJ0NdBziXRY1icpbgd8OwlIsJGWFX/sdeQ8NLe3mIc/1yE0iSZEkibV55OrDKZAX+XpDoVRn74+dc33fGid4rkdzbxTZoCXLsg13k3OcJwfZUkn0e30SHeckwTuat2pdo0zXGc9OB7SvDKbmsKUqsJ57Az9AFEZIkgRplh79WZ0OCi0agvNiscBkOrFi1Vrr9QJ1hAer5UGZ99EBx5phg+EAV1dXkIIEuF3PxeXlJeI4RlVWWC6XmE6nZ32ZeAD7vg/Xc5GmKQI/sHpTD85NbP/z/A+EJ3gWqdb1x+a3tMHNQUIIOIoCQmBNvO/C83sMLMgsJVlIVajW49H+cfi70w6YWYuPpUD20RB9ywDDLjggK7osy9Zdqkc+y20d1fbXWAx9O8PRpSBRCIE4jnF5eQmlqBs2CALa8PZ7MNpgNpvhx+0P1Nn5suTGGHge8UCjKMJiudjgy78bmLXN7Od8S2BlEaVIt9F1XQwGZL+aZRnynBIXx6z5nQ4KeRLK8gy3d7fwfR9pkq69fU+04LT15phLCHSXUySlhKMchGGIfr9P8gJparkYSimEQQghBOaLOYDzXYvWGr7vIwojWmDSFL7n70xxd9VakM+DtTA/0YJZu79wmaqsiMTehWf3GPh94MVdqrVDjeUTP5LN3vczeNNmF2QNO55eircad+1APkkSZNnDpqpD55JdXuy7pIvagWlXYkI+J8+lagw7vvD8Wlc1+v0+4l4McXv+ge/7PobDIQBguVjC9/wzn9F+4MrfJ8d3E22NXKUU4l6M/qCPVbLCfDG3G6tj0OmgEID1mE2SBHmW28Vmo4S1K+P0E6NdKs+zHLe3t5jP5/b7QRDg67evMDB20Tvn/RkMBhBSYD6fb57P1il1Wdx4ewE/9z3tCtr6mEoqaKNRlVWn9M8eA5cteYPJu2+ANjOHyIy0NxDtDmzXdSGEQIVGMqLDY4czd0YbVLra3IB397RfFdtJCNbQs9/H2gawC9lNz6Us4Xy2XhfegyLAJ56H67jQmjr3ry6vYIyhGGA2J23K6jjuZeeDQmDdCVrqcifXrwsv4VuiHVBlOXWTcZaQvy/FZvPJueD7PsIgRJqlyLJsrUwPdDqT9ImXg50StGnkhRqtrM4vQI1siBTk2uFImg4NDIQWqHV92NxiSC3BdmS3ZEwAoEK10/6vLZFz7rI7B4bb8+1Hm2stttacPM83xLcDP6DnK2AbAM4FYwxGFyPS+5tNSQuywbnH1SeOBxtAAMSHvr8nYwWWrDkW7yIoBEANIPphRpAn9N2/8rIXYJu42fXFbKOsuqO8JSXZSLGR+HPX85pBo5QkKbBarey5PJZF6vJ9l0rasndRFp8clwbMX2EPctabew9gD3Uekyxgz1/j7NA+gVA7eGJ+pVRyY25pZ2wsdaXdKLedQT9DIMbnI8zm9duM2YGvapff8aegjYYU0ioPbAt4G2PguA6SVXKWTXj7uQghsFwuybtam41n9YCi09HnwZsRxyU9yKqqrKXtR0dVU2f5Klnh7u4OeZ7bpr66qo/WyHw3QSHvWncN6FMQoIH3swuWStquXjYKb4M1i1jEmiezx/Ca180ZzKqq4HvUOs+luV3Zkq5CCom4FyPwA0ymk05rfb0VuHTMgWDbXairiw1DCAHlKCucXFc1yqpcu1Uc2cCmaw0ttPX45fdP1yQlsS2H06bAdMHOq31e2zAwkDhMOua9Zqq4OsPZ8O1udR7vaZaeJyjEWi+UG14A2pRHUUTUhbp6YGTQ9Xc1iiJcX19jNpudverVFUgpIZVEkReYTCZwXRe1rq06wLF4P0GhEFBCbex6dvHSPgLqukae55hMJiQ/kBcb3/cDnyav+jif0lOgLEooRZ7HzHHMctJTKqvSltS6PDExPM/DYDhAmqUbpaOPCgEqsXJm2vrBbjUPdPXZckZQa300D6cN7hDURkNirdNpXTta2cHHfv/c94y19/jv7crENtoNIec+79eCEOQMNZvOkKapFQnmYMwPqJGDhbnfGnZMsVxQE/vxu5nlGZIkeVcbcSEEwjDEYDD4nG9bkFKirmq4rguribklxv/Ue8jNZI/9zLsJCgGqn7O0gwEptNdmc5C3id4/I7hMoLW2DgDb1xr4gRUP3pDtOQOYvM+7vB8/fqw1FDvsN73L3tAYsmF6L+XRt4CjHPi+D8d1UBTFhiF7lyFAEjoQsO8JZ/WOPnZLKFhrDSWU3cCee5P2ErQXDOZFtuVitnUKHygG/IRobx7yIrcSOgzf9wFDgsvnmB/anfMbXzcG9/f3dkPS6blLPCxv67qVmW1BCvlhvcoFBDQ0hqMhHMextoAvCQj5+0Y8LhfWzRV5G4ICQschq7sgCDC+H9Ng2ZY0eSUZg+eO+2blHrMmgbdJ7Mz9iaIIvu9Tt3aeW27GOVHVlc0ktRtiPM97ekfTgXsexzGCIAAEBduu6yKOYgCwQdD2OPxoMDAIg9CKpnMpmQOtTnKYBHUEs5NGu3TLXMBjhpe9TrH+t1CUWd3epfPi1pV709blNDCIwgj9Xh+L5QJpkm7wIbfHvTan24Seu4S+jfZYbpfXgyDAaDTCKllhuVieLVjZHj98rttl166Ms21YmShHoRf3oByFfr9vdSDLsoQ2lAwpygK60u/iuk4NIQR8z8egT6oei/mCeNFVvXMu2XdtehdBIXc3sjZfHMfk8Zvn6x1Ew/15zS65LkxS9vo4BVyTxpoQAoEf4PLiEtpoIhqXx3ciHQsDyizsysK8JDNzznuulMLFxQW+fvtqZVeklFCOwnA0RFEUuLu9w2K5QFmWHzYwZJeXtsUd0JSyuulaBgC2U5qDV5bVgYCdYA99ptsNJW3xaiklYLq/iPH5e56HMApJZxTPOyZ0YZ58LWwHIZ7nYTQaAQAWi8VJaQjH4jE9yC7DcR1cXlzi67ev8DzPvjee5yGOYggpcHt7i9vb2w873wop4Ps+giBAWZV2jdVGn6Ti0fmgkJsqpKBJ23EduK4L13EtJ6jNp9jZzfeTwl6jJu2ifr+Pfr/Z0WeplUdgPbZP7AelFFzPRVWRO4wQazeTMAoRRzGW4RJpmm7IBHwk8ATFLjthEBKXtapR1VV3s6gGWCUrWw7lDKHrueQxWhze6dgOCFkaqq2JSB/fbW1V5hRy443rNvPtDpu7j5it0UZDSWUdTtI0xWq5sgH/Ry1tHgNOdDiuA11rLOYLUqpoxlyta8RxbMfiR92IC9EEhWGAelWj3+uTYUBZodY1six7snm2zSnc9b52OihkDiFPqNyoIBV133BJEmgmpgM7Bd89TNMEMRjAGIPFYoGqqsi6y1RUbv4gk/WpwJwzKSXSNMV4PN4QT7+4uMCXL1+sFuRHDAiBdbaE6R2+58PAWM4o85m6Bn5uAD1ru+l0iBt5TMOAMcZmHoF1gFDr99GdLUTD3W7+5CqNcmhzXuNjjvU22EpuNBwBBphOpuTjzJnyj7gOHQk77iBQVRVub2+xWq1skBj3YsRxDM/1Tsb/fa/wPM/SxH799VfUurYb8f/4v/9hf26XpBZzCh9Dp4NCRzn49ss39Ho965bgez4838Nvv/1G2kVZjsl0gul0agOhj5AlbENI8uAsyxLj8Riz2Qx1Xa81HLu7/nQXgjYhVVlBOcr6SgKUQWRiL3clfkS0AxspKHioK2qkCMMQRVF0NvhhvmpbWLrX70FKaTMQx5x7GK45lu3qxTaRvmtQSmE4GOLy6tJmY1zHJSrF6ALDwRB5nmM6nWI+n1sf548GIQTKkuwc2d3EZrU6/Hy7DCmJwyqkgOu6gKD3pyxLq7LBAs11VR+ll/mewRu15XIJ3yftXK6eKqUQhAGy9PCGv04HhcCad8bkyjAIqRtOSMshZB9AJrd/NNR1jclkgvl8jrIqrTg0d2b/rB2Brw0ppbUn4/HGt5IzApwVMvpjbUQYnutBQCBJEiRpAhhq4PB8r9OLYzs4E4JKVo5yUJTFSVwBqqqyHMJ2Y4YU0lrHdRGcreFOVs6gQqz1KCGoGcD1XJii22Xw14IUEnVdYzqdIs9zO2ZM/fHuxanAQXZVVjs3ZaxkUVbU4f0R51uAqGJxHKMoCiQraij1PA+Xl5dUSf2ZOYVVVeH79++QUsL3fSL0XpDFEFu78E7iFBP5e4QQ5LnJmnHMv6x196Uvug6tNfIi3/mitUWPpZSoRf0hS0ZcOs6LHHmeW2FVAJ2/HxzsSykR+AFlCYvyJFSAPMvXElot7s5jPJ6uoKoq3E/ukaQJlFKIogiXl5cASJh5MpmgyAu7+QQ+Do+wDSFJ8WG1WqEoCuvp/onDIcV6E75rPfcD4i4XRWGpGB8RcRwjCiP8+PEDd3d3pIcqJS4uLlCWxzc6dTooNDBW94kDHN/3LecnSRKbFbO8ww9WOmbbJUc5tnzHQtGfOA5FUeDu7s4KbrfBJWQWb+56WfCUYP6uAJV5WEy1693G2zDaQDjkbKKNps1lfXxjjDEGZVVajmLbe/Y9jBGtNdIkpWyg61Jwb4AsI591XWt7bazF+NHAAWBRFGj8aD4rMkeiqkkN4Pbu1krOaaPt5tJ1XQgpzqYFeU6wPJQxBmEUYrlcYjKdoKorRGGEoizIUvYEVoCdDgoFKAvm+z6UIu0imLVqe9uw/SO/j4EfUNOD0fjx44e162Jsc94+u5FfBqMN0oQkOMqKeGZBEFhZpDRNMZvN3sVCf2q4rovBYIAgDDCfz5GkCTzXgzYanushCAIsFotOT97GGMS9GIPBALrWmM6mJ3GkaGsdGm2Q57nlo/L3uyq+yyVi13URBAEuLi4QRqHVc+TyMrCeh5+aT7p4jafC6GKE0WiEm5sbJKuENoifc+vBcBSpiZQFZbu01jYL5vkeer0e8jx/NCj8WTO1VVVRY4nrI45jqxla1zWqqkKSJBhdjAA0pfX6uHeu20GhoA7QqqowGo0QRiGpyUvR6cXmraGNhuM6Vi+uzZX6xIFoaV4CxONgsd4oigDA7sp0rT/MpoQ72T3PQxRFMNrYUg83HTiu031va84+NM81zVJkaUbi0id8b7bFjrseJCm5nkNc17UC3wA2NuQfHVJK+J5P9ANB2qW6bIKYz8DwNGh6BzzPQxiGqKsaq2TVCf3dt4TjOFbmaDQaIc9zythrTbSFpjFHSEFBc0sr85D5ptNBoS2NOiRoWZUUFbuu+6GJptvwXI9KOZpkEsqitKK8XecwvRcISdmdMAgxHAyha207vDiQ+Aj3mTPzTN8oixJFXlg9Ps4SFkXRKSHfB2hckuq6xmq1wmq12ggIX/NZdjlosDJgUqLX68FogyzNEIbhZ5m0gRACnushjmMrkaYUZYbZdeMTx0MK4ifHUYx+vw9jDFbL1YfrH+ANZVEUWCUrAMBqtbINttyEK6VEskpenClky9xtdD4ohACurq4QBAG+33yn3avnbvo8ftA5igdLEASQQiIpEgRBQO37RWHtgD5xPIw2UK7CcDhEGIaYz+frjkOzth382cESPEmS2GYKAXLVgSGxedd1qZzWcZ9fIQSSNCEOYFl+iKD+pYijGIP+wC4+nB3vusbiW4AFlj3fI8kqRdxLJZXldbW7zj9xGKSUcB0Xvu8jCiMsl8sPGXTXdQ0lFcqyxB9//IEojGwvhVLKWnYKiA2ayq771JbHegydDgoBKu8M+gPkRY4sy8h4HDRg6rr+kCKWbXFc1lhTSuHy4pLKGDVlUZeLJf744w9SOP+coI6C53n4+vUrvnz5gvlijvF4jCzLPtwYZGHejW7LRjTecRxcXl5CCIEs3+0J3bVxyKWoLmfv3hLGGHguWbfVmrKoURzZDCKAD58t5HKdFKSK8csvv1g+bVmW+P0fv2OxXJz7NN89XJdcugaDAaqqemht+0EgBAlQOw6Fa3mRWw3isizxt7/9DXEvxv39/YuSQBsJtR3o7EyojYZUElfXV3BchxooytJyldjyzqDx/DMfs5zsueRLqhwFA2M1xpSkBh3Xcz9U0PJaqKoKSZrgfnKPHzc/MF/MN0SOuxbsvBYMms7jVpnVyroEAVzHRZZlKPKi87zftwwE28Exz1ddhJQSg8GA/OXnc2Q5bXx0reE4pOX4CSAIAuvN67keyooEluM4piD6g8wHr4k0S5HnOeq6xvh+jMWcvKW7+u68Jtrc5HaTWhRF6PV6KIoCi+XClo4fyxKyraedj3YM05O/4ceWizTWF2MM8VkmmoSZe70eAj9AVVfrDqT2x5nTnMM5sM8kYn/WAJ5PdjdZmuFufIe6qhGGIa6vrwFgQ84HeDql/NGwzz3XWmM+myNJEmtr1w4GH7uHj33Ge77n7WvijJFU0lIXlqslirLYeY3nvO59nvepvYl5Im+XX7s2BoSgBr5VsgLGJEHjuZ4Nej5i6W4XuNEqyzLc3NyQNpwArq+vMRgMbPfsJ46DkjSX5AWVRHfJRXXtHXptGEM0prog95x+v48wDLFYLCwv2orPvwDvilPIdjbfb77D9304ykEYhvB9H4vlAlmWoSzLjSzYR/H4FfyfJIKp0QbL5RKr5QoQ1PgQ92JIIa010Ee4L6fErhJZVVVWFPwjZQefg5ACYRBCCIE0pd39sbIIbw1t9CYv9MRrTTuY6vJCpmuNyWSCxXwBP/BxeXmJIAiIvpN+PLoEoy19xtqNy9XSclLzPMegT9JGVf2xGiFeC+znWxYlhPyca9sQQsB1XERxhCzLMJ/PrZj8sxWahu7zGPYOCl9rQns0q9DIIDiBgyzNcFvdIkkS0jBs/JDf4vy6BCGJYOp6RMItyxKrZEXdnoZ0C13XRZEXcF13Z8r9I9yn5/DcPWhnrduWd1mWWTmA9nF2Bd8/431uX5MRxvoGB36AyWSCJEk6uTBuPwuNTfkQGxg+8vPHfCbv3g/NFL7FBoQb+xzHITu+skKRU5f5crW0jklGmw/RVLUNAwPXcfHlyxcEYYA//viDyptVDdcj+Z6qqsjzG4dvGo81YHisq/Q9fHZ7ndJaw/M8+95AbM61P+Pcugu7sqNRFGE4oKbH8Xj8oPHxuWPZIPstysfH4sEFNZ6bRV4gyzKrDWfJki1+U/t3f/YsjlQScRzD8z0kSYIszawkiOu60LW2Qp8f5eV5TXheQ76vyYg9L/KdO7KPlpV1XZc6soMQSZpgtVq9mzFnjLGBoeusNfnY3/cUdnftz3pJ518XoLWGETSOJ9MJptOpFRK2eOEldP1aXwou/3NT32q5Qp7lVqPU8zwoRyHNSOyeqQKH4pjfPXb+eevPfux3XMclP19HYTqZbnTWfmRorTHoDxD3Ysxnc8xmM+u4xRSQY8ZA5ziFu4SXq3pdtmvvtp/a0byXyWg7oH3Jw9Ra2zJOURSYTZtBwZIgnou6rkk2pOFjbH/Oe7k/r4l9XhxHOYijGHmeYymWtEhs8V/tuHzB5uQ93//2NTmOQ/yqPMP9+B5Znr1op3oO7HoWHBgGboCv377i5uYGq9Xq5J/dDgq7yikEHmZgrIVoU3J6jmv5IFP+k3SK1qhtFrUqKyyXSzvncsXGcRwsFtR1vM3l3hcfJSgUEHYDsn0c16PyKFOldq33XXyHXh3NOq9rjcl0shEs71qD9oUD0C6oNOtOSq016Y/p1xdy3cZjC+pGs0TzwvFgec+ZmUOCQv75xXyBpVgiSRJoreEox2rDlVWJoixsZms7TfwhX6YtPHav2/drQ8y44WvWdf0o4f7BfX3kNr/XTnmecPi+ZFmGyWQCgIR73+NltctWjnKsp+9jmcJ9giL7OxwciePfvQcyPyfSyLSdidgsc3PWq/11WyIUO8jqO67xvY53C0OND3VdYzafEUWirOA4DnSt4TouyrJEmqTk2Xskp/aoMXLkWHjLz7ZqBs0Y5j+NMZaew01rH8lf/iloo7FcLpGsEqyWq/3eLbN+F9tJtramLGUKm10gE8Z7vZ6tOT/Gkdq32/ITT+Mlg32j61MI68AQhqHdxTqOA9chx5cgCABDDRLtgfMReG8vwWNjlTWgeMNh77Gh34mj2N5TnqjaCyoAevmeCh7eKXHaTt7tDVvDMfMDHz78J3+/a5lCgK7JdSm7HkYhhBQ7NRYtWl9+kPVrfUQ7cOLf4efepr88i9ZELiAeNEG9asDVOm9utmjzznZleIDdPKj3Dr7nVVXZrmygyWq5LlarldUwPFa655h19Nh73ZXPDvzANlT0ej3LL2R0XRz/NVGW1OEeRuHLf6n1LtsAsIkZypI8k6WUFBRyFB74AeksRdFGBu5Bxs48PhF9FGeHU2Pvwc0/zuo0xsBRxHfRRsNo8i4d9AcPfvUzKCTsnPzEjoUOjW9tQ3z2XO/xMc4x4TOE7Xcrltzazdt5gIObVpDTxbL5U4udFNI2EsRx/Ogcx2Nh4zq3NwCi9bMtRYQHgdwBQSH/247TRz77ZGgtJFKsm2XaQepGINxkEX+2xrbtTBaAdbWqFQjzRvxnCczO+dlaU+OXchUGg4F9f/hnNjZunzHHiyDF2pIRgJ3LrHWgaTKFPHmVZWnFItm+amdWAI8//M9M4WHY92VqLxJaa+qGlYpErDlrZYydzNsyEp9BIeGpsWpgNvhQxhjUut74Ny8KvFhwiZm/f+hndxkbiyN9wcJmv/D4prGLQSE/O+Yp83y461w5KNxYjEzr2M9sFrYDqJeCx9pBn30CcPac34vHMoW82dneFP0sc8yupAe/C7wB2BUU7/sZx8wPP8Nn8/vHTRO75punklOfeARbGxbmbtY1cWYhOChs8YOyLENZlRs6bNs73CfLYkdmCn+WyWNfHEtK5myvtaLSa54Ucy8/sYntbN32ImazQoDdHPF93eBWtbJGuziiO4OLdxoU7sJLGmt2/exb46nnzc+Sgx5ttoTx7Q9u/ZOzdTBP/vyDRW0vGtDurOKzn30C7Az+zCNfb/97e3Pwzqf1bT7ldiWtvZHYCJo/U1gvwoP7tV2xaTY/Usr1fW79v/G7Hwx7B8atH5dSIjCBNWOQolU+llKuG0yaxe2QEtcxOkXApjbcJ16GXWKyQglIrHftT+FnClD2wfb4bu9yOTMCbG2EJKCgHtyz7UYh/rNtSbRP8PRe0G5IAJ6/rnNe91PPG2gtTFJAQb08gBXPL0iv1hH6gs8+Fg8+u/WZj2UK7e8+k0R4T3iqCbIdJAu1/t4ha+ix9+wYaso5PvslHe3tMf6AlrGD5vbRcOgzk1JCSQUpqZoohMD/DxGQMKjLvlROAAAAAElFTkSuQmCC"/>
</defs>
</svg>
